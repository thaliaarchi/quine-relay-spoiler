module QR;initial begin $write("%s",("let s=(\"Module QR\\n\")\nput=s\nprint\nlet s=(\"Sub Main()\\n\")\nput=s\nprint\nlet s=(\"Dim c,n:Dim s As Object=System.Console.OpenStandardOutput():Dim t()As Short={26,34,86,127,148,158,200}:For Each d in\\\"BasmCBBBCRE`F<<<<C<`C<B`BBD#CXwasi_snapshot_preview1Jfd_writeBBEEDCDGECB@IUDHmemoryDBH_startBDL|DRBAC BAJlACA4RB9MiCD<AERCA>D!BE@ABRCABRCABRCAJ!CE@ B-BB CACk:CvACqRC COBMADRCACRCADRCABRCABRC BACj:B-BBOBMADRCADRCADRCAFRCMM}CBABM~(BBBCBBB,BBBDBBB0BBBDBBB4BBB=BBB?BBB;BBB ...\\\\t..\\\\n..(module(import :wasi_snapshot_preview1: :fd_write: (func(param i32 i32 i32 i32)(result i32)))(memory(export :memory:)(data :\\\\08\\\\00\\\\00\\\\00$:))(func(export :_start:)i32.const 1 i32.const 0 i32.const 1 i32.const 0 call 0 drop))\\\":c=Asc(d):If c=36:For c=0To 11:s.WriteByte(If(c Mod 3,Asc(6"));
$write("%s",("24163.ToString(\\\"x8\\\")(1Xor 7-c*2\\\\3)),92)):Next:Else:n=(c>124)*(8*c-40304):Do While n>127:s.WriteByte(128+(127And n)):n\\\\=128:Loop:s.WriteByte(If(c<125,If((c-1)\\\\7-8,c+66*(c>65And c<91),t(c-57)),n)):End If:Next:For Each c in\\\"<?xml version='1.0'?><?xml-stylesheet type='text/xsl'href='QR.xslt'?><xsl:stylesheet version='1.0' xmlns:xsl='http://www.w3.org/1999/XSL/Transform'><xsl:output method='text'/><xsl:template match='/'><![CDATA[sub f(s$,n)print(s$);:for i=1to n print(\\\"\\\"\\\\\\\\\\\"\\\");:next:end sub:f(\\\"\\\"write,format=\\\\\\\"\\\"%s%s%s%s\\\\\\\"\\\",\\\\n(\\\\\\\"\\\"\\\"\\\",2):f(\\\"\\\"write{-}{txt}{echo -E $'(\\\"\\\",1):f(\\\"\\\"\\\\\\\"\\\"with Ada.Text_Io;procedure qr is begin Ada.Text_Io.Put(\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans B(Buffer)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f("));
$write("%s",("\\\"\\\"\\\\\\\"\\\"trans O(n)\\\"\\\",2):f(\\\"\\\"{\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"B:add(Byte(+ 128 n))\\\"\\\",2):f(\\\"\\\"}\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans f(v n)\\\"\\\",2):f(\\\"\\\"{\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"O(+(/ n 64)107)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"O(n:mod 64)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"O v\\\"\\\",2):f(\\\"\\\"}\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans D(n)\\\"\\\",2):f(\\\"\\\"{if(< n 4)\\\"\\\",2):f(\\\"\\\"{f(+(* 6 n)9)48\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{if(n:odd-p)\\\"\\\",2):f(\\\"\\\"{D(- n 3)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9"));
$write("%s",("):f(\\\"\\\"\\\\\\\"\\\"f 27 48\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 36 11\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{D(/ n 2)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 21 48\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 48 20\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans S(Buffer\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"STRINGz:=REPR226+REPR153,a:=z+REPR166,b:=a+\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"2\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"+z+REPR160,c:=b+\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"8\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"+z+REPR165,t:=\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"class QR\\\"\\\",2"));
$write("%s",("):f(\\\"\\\"{public static void main(String[]a)\\\"\\\",2):f(\\\"\\\"{a=(\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"write(\\\"\\\",4):f(\\\"\\\"'implement main0()=print(^1^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"BEGIN\\\"\\\",2):f(\\\"\\\"{print(^3^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"echo ^1^\\\"\\\",4):f(\\\"\\\"'f(s)\\\"\\\",2):f(\\\"\\\"{System.out.print(s);\\\"\\\",2):f(\\\"\\\"}s=^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"389**6+44*6+00p45*,^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";for(c:(^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"#include<stdio.h>^8^"));
$write("%s",("nchar*p=(^15^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"Ra#include<iostream>^16^nint main()\\\"\\\",2):f(\\\"\\\"{std::cout<<(^31^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"class Program\\\"\\\",2):f(\\\"\\\"{public static void M83abbSystem.Console.Write(^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"Quine Relay Coffee.^64^n^64^nIngredients.^64^n^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");for(int i=9;i++<126;)[3pva$^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",2):f(\\\"\\\"{i\\\"\\\",2):f(\\\"\\\"} g caffeine \\\"\\\",2):f(\\\"\\\"{i\\\"\\\",2):f(\\\"\\\"}I3b54rja^64^nMethodv4f#aeach(char c in(^6"));
$write("%s",("3^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")))^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^32^[2al3dp3c[2cs3c,3l[2k@3kqa^31^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")s rts(ecalper.h3eja^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"     53c4a SUTATS(egassem^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"rts(nltnirp(])]^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\".NUR POTSu4cba.C3dh3dX3bba[65bX4df5lp3lna\\\"\\\",2):f(\\\"\\\"})1(f\\\"\\\",2"));
$write("%s",("):f(\\\"\\\"{#\\\"\\\",2):f(\\\"\\\"};)06xt3dba;+3nna3(f\\\"\\\",2):f(\\\"\\\"{#qp]^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'[p]#3sv3r23)ga7(f\\\"\\\",2):f(\\\"\\\"{#.33)ca51h4-ba1S4w23F?7d33&r7u53sda,4353.ma^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\"));
$write("%s",("\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"' D ; EYB RCL4/v4+ja36(f\\\"\\\",2):f(\\\"\\\"{#DNEm4[m4ada. A~5[p4deaPOTSn4[#5e~5[o4boaRQ margorp dnex4[x4abaS*5[m4c2<[ca91j4[j4eba&%6[l4bgaS POOL)<[:7dba^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'j4[j4[j4gda&,)(6[?>cga. TNUO<7[s4bfa(rahcg:[(5dgaB OD 0B>[t4cca&,,<[,<aca)A36[;=e6=[.6cqaEUNITNOC      01z4[c9c,5[W8dK7[aGeeaRC .p4[p4aka,1=I 01 ODt4[TKecaPUq4[/I[6<hva;TIUQ;)s(maertSesolC;^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\"));
$write("%s",("\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'Ye%4Rra744(f\\\"\\\",2):f(\\\"\\\"{#tiuqn\\\"\\\",2):f(\\\"\\\"})215>5[qa^32^\\\"\\\",2):f(\\\"\\\"})959(f\\\"\\\",2):f(\\\"\\\"{#n\\\"\\\",2):f(\\\"\\\"})420pY4d8,ba8AAbg8[da304zY[O7bda218lK[wL[j4ldamif+6[ga)91361\\\"\\\",2):f(\\\"\\\"}5[,6[j4lbat(6[(6c%a315133A71/129@31916G21661421553/04[04cva%%%%\\\"\\\",2):f(\\\"\\\"}*+1%%%%811 -\\\"\\\",2):f(\\\"\\\"})48\\\"\\\",2):f(\\\"\\\"{3bhaj:+1 j@34[34cbawm4[m4cl4[l4cbaWm4[m4cba\\\"\\\",2):f(\\\"\\\"{m4[m4cva)(esolc.z;)][etyb sa)t=[#>[j4[<6hea3289m4[x5[j4lba,l4[w5[j4hla!\\\"\\\",2):f(\\\"\\\"})46(f\\\"\\\",2):f(\\\"\\\"{#~~v4[%5[j4hea(rt.o4[z5[j4hba)A7dda\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"};l3efa~~dneo3hra~~~~PUEVIGESAELPnr3ala~~1,TUODAERw3a63j$a(etirw;\\\"\\\",2):f(\\\"\\\"};u=:c;))652%%%%)u-c((||13jda#-<q3jda||i)3mhaBUS1,ODs4qka)3/4%%%%i(N4cx5kU4xPa2=:/t"));
$write("%s",(";2%%%%t+2*u=:u\\\"\\\",2):f(\\\"\\\"{od7 ot0 yreve;i-=:u;1=:+i\\\"\\\",2):f(\\\"\\\"{od))1(evom(dro=:t elihw?s;)s*45oi5vv3jd7dladohtem dne.s3dganrutern3d~aV);gnirtS/gnal/avajL(nltnirp/rZa|atnirP/oi/avaj lautrivekovniJ3d.4j[2cib\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"};0=q;)]q[c=z(tnirp.tuo.metsyS;)0(tArahc.y+z=]++n[c;y:]q[c?n<q=y\\\"\\\",2):f(\\\"\\\"{)0>2%%%%++i(fi;48%%%%)31-)i>3c&as(+87*q=q\\\"\\\",2):f(\\\"\\\"{);82122<i;(rof;n)rahc(+K4r[2k*3&oa=]n[c);621<n++r4aqa0=q,0=n,0=i tni;N3&bc6ayi4asdRbQeslxfvfllRf<bedRb;fr6;agb-a|dzdxdRfGb8aqeRdYd5aDUGi;agb-epb>aqeRdHa>aJaRaAdteFbaeIfOa5aac2gAz6f9azb<a4aLa7a;a4a<aPhsmkdxd;aNa?c6a|eebHaFaIaebzeJaeb9a/a6a2dQbUe-f2a-I3bga5d6cRbE3gdd-f/aof0fRfhpEkEf.b2e6aRa;dNaxbogO*Gh;aTapc4aLcEeyiof6amc<byg-fJlsbvh|b*bWfybxcxc>aGaUeAa2a6a\\\"\\"));
$write("%s",("\",2):f(\\\"\\\"}g7a6a@a\\\"\\\",2):f(\\\"\\\"{g:a?aMbKaKa6a?e:a@aEa2a|gZfMbbgli>a:b1a-gqmUf\\\"\\\",2):f(\\\"\\\"{bHauc6.0301O;01EcB6JaMa\\\"\\\",2):f(\\\"\\\"}bJaPyEc-bJaJaUa-bJaMdJa8bTr;a8bjuKa8bjucWwbDWPaOaXtNa+b9bKa8bSaNa|08b9sju8bNa+bf4JaLaJa8b9sNap4c\\\"\\\",2):f(\\\"\\\"{3aia03+b:bO;.4agaDWJaHa\\\"\\\",2):f(\\\"\\\"{3ccaf4m3a+aFdf+;a8bSaUa:aUa:aTrviSfQfRl4aM/sbsb2be3^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'oaviDa-a|b*b*b-aJ6aua?aGaUe>a5j\\\"\\\",2):f(\\\"\\\"{gKaKa|gZf,6cgaagQjkg06esasbvh*b-a/bxcHa|fNke3c2c\\\"\\\",2):f(\\\"\\\"}b\\\"\\\",2):f(\\\"\\\"{gph\\\"\\\",2):f(\\\"\\\"{gvg1a-g\\\"\\\",2):f(\\\"\\\"{bHaNkRf-e:a:a\\\"\\\",2):f(\\\"\\\"}bHa?a\\\"\\\",2):f(\\"));
$write("%s",("\"\\\"{gJa\\\"\\\",2):f(\\\"\\\"}b5aAdte@a1a-g0iNkxcpb7anb2b:b\\\"\\\",2):f(\\\"\\\"{g2f@j@d-aIfekxcHalgjghgmk-aUf0ixiRf-f-gSf|fNkzeSgxiHack;a/aDh<b+hWh<apb/aDhWhnb<a<a7b:b\\\"\\\",2):f(\\\"\\\"{g/aDh-f-g+gFa,i|b1ali3b:b\\\"\\\",2):f(\\\"\\\"{g9hHaNkHaUe-iCe|bxc3b0a:b\\\"\\\",2):f(\\\"\\\"{gIa|bzeJa|e5buaQbxi<b=a-aHm*c3bxdUem3aea|b9ai3eta2bMa7arh|bphnhlhjh9m3hAaAd7RPcgfvfOhJh7aEa|b8k6kMaHm*cEc,dJa>a2aIfzjMgMaHm|b<i+cbi6a13kYaxd?Bvb8g/aDh=apiRa-*Cd-*0EN9,hDhsk6a7b5ackRfwb\\\"\\\",2):f(\\\"\\\"}jUe2b5a9gYi4b-bhc+sOiOikv0c/bxd;a<hoj=?aea6a2bi?eucQDDR6a5n2a5awnbM\\\"\\\",2):f(\\\"\\\"}gEhglCtOi6aUhvnHa1dmdLhRfXkJkHa:eXkJk;l<b3bxd6aIhDkPh4lU/kixb9iacPa;aXiccq\\\"\\\",2):f(\\\"\\\"{pbub|bd+ZboVnbpgujsjEc,d?aRiWkuhUk4j<b<b<bFj:b<j<b<b,cKjHj7b-bKj8vSg3bDd0kMi9a7b6g-a5bM5,cKj=a9a7bubxbs3e33ecaCj33cear=8fC3c13ifaJb7bdU3fmab8Eamh9a"));
$write("%s",("7bH2u3amakiykpjCk,cKji3asapmhh.bfh,cKjsbHa\\\"\\\",2):f(\\\"\\\"}g\\\"\\\",2):f(\\\"\\\"{5c^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'aVjDjCaLi6aakflhk4j6aKk8jYjel.k<bzefDc93gca;k53cIaIkGk3a6a<bkicjaM2b2a2aWJekZk0iwb\\\"\\\",2):f(\\\"\\\"}jRf@a>anc:e7b5aWf=anbekyb\\\"\\\",2):f(\\\"\\\"}k5a,bJa6awAa%aub9h5aUgwb\\\"\\\",2):f(\\\"\\\"}jHa:e-b9a9b9apkekyg>am3aya5Jekyg@a>a:a|b9a0b9a@a>aaCaYa>e|bPg9bJa0bekyg-b9apk9aCaAaJa9beknbJa6a|b5a,bRf:e-b8ka|-ajh9apbkvRB9XviWJyg8bAdGh-as3anaSH.bbb-aWJyg7y3n5aWJKc>iwXxd6a-b9a8b9a7bJcJayb>a8Ski>aJa*c@dxc?b\\\"\\\",2):f(\\\"\\\"}uo3a3a-bIlteUe@a>a<a2b5aDcd3:atcJaub5aEcd3?a,b4b-bVgs;aiaTkRkmdLh77"));
$write("%s",("gwcdlblpb;awb\\\"\\\",2):f(\\\"\\\"}j*l\\\"\\\",2):f(\\\"\\\"{iGTDR4ZERAV5ZH@3ZJdHd,l2nInClmm9n7n0n\\\"\\\",2):f(\\\"\\\"{vInVly>46IrN+Gu:rR5CL0xabbswH3xwH\\\"\\\",2):f(\\\"\\\"}brK\\\"\\\",2):f(\\\"\\\"}Mc-qywUG6@WRC7+RNn:1zUn/*h.TFUn-73bjbAotrUx-tCa<yd5<5=aDahbgol5W<y>dG\\\"\\\",2):f(\\\"\\\"{LstAaYaHkDaib@afbh09b=@YpM/0pvujb=lX4cud3UKpS*v.9bn<<yJy>Dm.iV|7N1,oT|=a=6-Xvbkbm5YptbmbTatHOakqTaeIJ|\\\"\\\",2):f(\\\"\\\"}2WS:vkxsv0wd;E+bpA@1zuyP1bpEzG9,3/b29kBjVmbTa2qjb>o+bUiYax8S?JytqM8jr>tb.uwKLhc\\\"\\\",2):f(\\\"\\\"}vr=OjX+iP?Wjbdb@xrg\\\"\\\",2):f(\\\"\\\"}7?afb8ql+CCK,.0??nR1KS*ib+bkqhc3t<xjbHt*=zbAa0v<8?aw=zb@0r|eZX+AzValuPyo3y1db4b<Lh|?EmuzZ-jRNZaG51v2p\\\"\\\",2):f(\\\"\\\"{xp5|bLxK:eOAE*ba~6fxdDa1Kvqzb454ICtd5puh.ykrR<aNz6JG9E8wTmbG-4bQa5Hs68usyUxrmbbyolu@LGubqG+jsyPVvh9<z/bZEjb0z1pWaMEbPjS3bMy5bhbe95b\\\"\\\",2):f(\\\"\\\"}b?qqy7v.9g"));
$write("%s",(":tbk1O/j66b.vYa\\\"\\\",2):f(\\\"\\\"{;O@,b/@Raf@zvub.bQzlblWac;pooIpgbWWx2\\\"\\\",2):f(\\\"\\\"}bytstAaMoH8E\\\"\\\",2):f(\\\"\\\"}hbCaMo.E03s>ZnD|W1wHvbeKJvT,kiCySaS?.b2rzUSa46EzqFDajbzEX7+2w76WwOc?W1wHMxXaFafrwq\\\"\\\",2):f(\\\"\\\"{+a?ykwH>o\\\"\\\",2):f(\\\"\\\"}vT?$6evbO+a;1yi;|oVaAa=4PpTaQX:T3,I>;ZGSy8S?2Vuw@9a?M60bOVj||oAamQv8\\\"\\\",2):f(\\\"\\\"{ocKC\\\"\\\",2):f(\\\"\\\"{Na5\\\"\\\",2):f(\\\"\\\"}3\\\"\\\",2):f(\\\"\\\"}1\\\"\\\",2):f(\\\"\\\"}vbiov8wH-twHL7vx9bEaz1jbFmgbCqCaNaq3aTb|rN-ZE8n4Tq5VamombNawHL=jbAo9v6Xv4UaFaPAmomb.b51ZEjbPycA\\\"\\\",2):f(\\\"\\\"{xNawH|G;O<?@0-bWWzUebkQy85>ZE46vGio?UwHxjlt=8ILM+jbj=jukiW@WW?H.b@W<Sjuc|x:<yvbioxbEUdKwH,wUaa\\\"\\\",2):f(\\\"\\\"}orCwB,Pa2Vv|sJa5adaLR2K9fLb7bubDa7blp<yDa|o7bx:<yDajr9MRwsJubir=tgbCa3bh@R9?afb9b6LZ6\\\"\\\",2):f(\\\"\\\"}brgxb2js6W>60=aRshbc>wR0bCaoRCaDah,S2x>?aDa<J;O2be=zWhs7bM\\\"\\\",2"));
$write("%s",("):f(\\\"\\\"}wAJAAslqpy8o6o<a,b4b<JTr@EDa+QNaY;X+1p;km3a\\\"\\\",2):f(\\\"\\\"}aDa<JlYS\\\"\\\",2):f(\\\"\\\"}wAdlDa-b<ajbebM+hshb^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'3crbn/eqV8yhDajsYao\\\"\\\",2):f(\\\"\\\"}mT5zz6.zdloI-GDa+Q\\\"\\\",2):f(\\\"\\\"}QT60*43v:7bibZp0?ZaFaNayEVPgbs61\\\"\\\",2):f(\\\"\\\"},p\\\"\\\",2):f(\\\"\\\"}FzUebNY4bEavy5H+b4\\\"\\\",2):f(\\\"\\\"}T@rm2qhpfpm\\\"\\\",2):f(\\\"\\\"{PX86eOcNaxbOp5V1HY<F1x\\\"\\\",2):f(\\\"\\\"{4ShbdG2R?a1pmb\\\"\\\",2):f(\\\"\\\"{bp\\\"\\\",2):f(\\\"\\\"}XopsvbkLDa=T7U/O@4=7Aw\\\"\\\",2):f(\\\"\\\"{o\\\"\\\",2):f(\\\"\\\"{/Fzi@Damb\\\"\\\",2):f(\\\"\\\"{bixQ@YaNwWz<B;kRpxh<B;kDax\\\"\\\",2):f(\\\"\\\"{kqhbRaeoubWSR2sRcl51.S<=NrfzhbKq|b?L5sWa"));
$write("%s",("bS2R?a3RzRQELwiD|-A*v6ub<G3oQ@*3X,mE0+ubDIrFpo/U/4kx6bv|ixjbO2-bY9<0\\\"\\\",2):f(\\\"\\\"{LrmFaOCqNHpB;L5@L/b|b.u,bksBMPaW*oJL|mW>R>7$Fa+aw|3,+q;2vb?aGa+U58>p=tF4k+NaxbDa4tibcW,6exdYa?.tb-vazb>y@Ta|B8UM6e5i;jbxxM4X:oQFaOvTEJOl=lbVzdrab2B|:apZXAfO@kG*3Aa5vpyjpubfN@Zs+Oa+\\\"\\\",2):f(\\\"\\\"}IY8|NVvv<-Tajptbhz=qUvab\\\"\\\",2):f(\\\"\\\"}B+HGaPHYu1kHpMzcvwtnpKx8|uZBaAoybjbaba\\\"\\\",2):f(\\\"\\\"}L/Ao>K.VHOUGybpF4|YabAu=ydPZu?D+FuNrdzhX1hhb5bH.IYOVDy8+SaP/OaEj||;*,b6>yru;/bZRYar9rAO=Ua|Wzb|WGVUGybzb4bRq|bEs3Jr\\\"\\\",2):f(\\\"\\\"}7+HdHsQndWmw3/$6e=gS*VsIAGtbtk\\\"\\\",2):f(\\\"\\\"}yd>G=+?=hsasCavb=32|uwMstt>,*rU*4U2UUaBfCa7=K1\\\"\\\",2):f(\\\"\\\"}|.bY|L+TazbXa;ObbFuwbGaT/evT*2Hm0U5D|RSkiO=M=qxVa\\\"\\\",2):f(\\\"\\\"}r=1Ao9bnoUtt7.8AoVUWalbHK0bNwcX,.>R|z\\\"\\\",2):f(\\\"\\\"{bDA1-+QQ\\\"\\\",2):f(\\\"\\\"{:T7F6b9bhbdbMo9b?a;A"));
$write("%s",("L|qJ7qQ=SCO=M=er?aArG*v;4vwb<?vb7kbv6sBvZoWaB6tbL2ZlZ3ybEaaHj,tLyZV6zW+/An>,O8bm5bAwR5g7m3-/Rzk+1hT9Ar<aXyBVTDCRp8RB9Xn8@z0b8yb-JA5YMr+77v9-yth>vx+bPSZ*z\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}bF\\\"\\\",2):f(\\\"\\\"{J|JAGa9*CaRSfV\\\"\\\",2):f(\\\"\\\"{AUwh?DI\\\"\\\",2):f(\\\"\\\"{x/pAo/b*bgpzb5W?We+p\\\"\\\",2):f(\\\"\\\"{=FxumdHKw7vT\\\\\\\"\\\"),\\\\n(\\\\\\\"\\\"bbnFm;35;AtbMxeEM><a5\\\"\\\",2):f(\\\"\\\"}3\\\"\\\",2):f(\\\"\\\"}Y|0bCatb0bxh?|T*Dp58c2D,,*UwWacbHpRSPpkiCyo?xsg:,bF\\\"\\\",2):f(\\\"\\\"{UXvt2bvv1|fx*4;+Tq>5;ZSaFuu1|75xoS1khqTuPnvbibN7|b6oD0:8,bp=/y|-y6G9Pa1|Faub|SMxB,M\\\"\\\",2):f(\\\"\\\"}K\\\"\\\",2):f(\\\"\\\"}6bj\\\"\\\",2):f(\\\"\\\"}D?=a24vvfxd>6pdy4b.MJ:E9epdmzK+A\\\"\\\",2):f(\\\"\\\"}GymzK+a54+7kPPp19=7qrBhT,7T*33<a+2d;fRDaNaAoPayk,|bP?aPvyIn\\\"\\\",2):f(\\\"\\\"{jwibWak.-vK+a5UaMyXaS=4bXaSa4b2j-37k?|.bIvRaUxp+2?Jv4bXaUET*<p\\\"\\\",2):f(\\\"\\\"}o"));
$write("%s",("Fajpg:kb8ye0dbjTy@7=\\\"\\\",2):f(\\\"\\\"}Bt\\\"\\\",2):f(\\\"\\\"}Ea+bbGatt2r2Kso2h,p\\\"\\\",2):f(\\\"\\\"}g4dG/bluT|czub|bw5cb<Y>,M6bS/bT@Wa9gk\\\"\\\",2):f(\\\"\\\"}Ny;p:tpsvb-BnZJ,FajtP*/b|b.yHV@Gk\\\"\\\",2):f(\\\"\\\"}abGa<SwbbSe|ltn|yb<p==c|cz?ajsd6aga2jp+k+(6epdgCtuNaxbNaV;W@2bM,CV?S>oAo3RxrF<\\\"\\\",2):f(\\\"\\\"{/Wa|byLw=ZaVzVttbqQC>zZ4bI,Eaft3,\\\"\\\",2):f(\\\"\\\"{4R3kb7rWaw4R3kb0I.I+QIy|bxusm,*WL+Hc|Qa<=fbybSY|4px-*1kVajuw|oVbo3besc2hb<6xuBvaB0RLX|b1zfP9bRa\\\"\\\",2):f(\\\"\\\"}*+;u1+xH|Y<\\\"\\\",2):f(\\\"\\\"}vu|\\\"\\\",2):f(\\\"\\\"{,VZtbjw?7F2J|dlWDcbwRwb9b4+8R2*7|Na>*Gp*bzbcr,bcbDak.Daaicbab49FgL<ICK+a;qxtu=62YY/O54bX7G5a;fbAou3alaXag2SazbdbjYQhxdhbd1pzo0;-PaqNPaOa=7z6/NrgqurgY1vYfRo0M5wJaiPP?4tbpUPP|fYrp1A6\\\"\\\",2):f(\\\"\\\"{6,K<\\\"\\\",2):f(\\\"\\\"{?HfR=WDzkC\\\"\\\",2):f(\\\"\\\"{|dbo5ybaZ0bebabPa+=z<juiDFaSyorwbI*Ns=.HwGa9*"));
$write("%s",("<0hb\\\"\\\",2):f(\\\"\\\"}JQaw4?@<aXyvb6AFaY3lt2bRaors7kbMS56xChbK/ybp1<04yu\\\"\\\",2):f(\\\"\\\"}LhJ|o@O|\\\"\\\",2):f(\\\"\\\"}oXar=Wabbe\\\"\\\",2):f(\\\"\\\"{mbK.TEk23bh<?.=F=4Cuq.z+hb7bB->tS4Ba@sy64J.VUVib\\\"\\\",2):f(\\\"\\\"}o**J9ujG97gE97bKLDE0vnxYZgP<a/0QrF;$6eOc*4=yKyhRV3x94uN5ORI0Xa??ro<0@CAaZoWaZaW:BvNZZaXw9bFzDzki9C+btLXwp\\\"\\\",2):f(\\\"\\\"{GFzb3br|U:8+ibuj2Hl\\\"\\\",2):f(\\\"\\\"};Atb-o+X/U<6mbwvstlbr|8:dW\\\"\\\",2):f(\\\"\\\"}u-7KXgs2B+rYq1by<7bibvt\\\"\\\",2):f(\\\"\\\"}b3hiNK5\\\"\\\",2):f(\\\"\\\"{bOabb*=dz8UWiPrj0+XDUFYxx\\\"\\\",2):f(\\\"\\\"{ZCL*=\\\"\\\",2):f(\\\"\\\"}bNaFYr|K/Qanyd;8UCL6qQsV;yq4b44Qag7rrFazb?yU=QaDakr3b<a*wubzWPaAoybvbbSe3a*a,*s|2blQt2bSRnIvOvboZaubJq19f;OvQ1Y3j#=fjbeK?aGIkS<pYsubIJ\\\"\\\",2):f(\\\"\\\"{6\\\"\\\",2):f(\\\"\\\"}vWalpP.|bKo5?8blbssBCHO*-ab\\\"\\\",2):f(\\\"\\\"}k2hkbnZr.yWJq=aJr,SXap/p.HOwxs/>i\\\"\\\",2):f(\\\"\\\"}"));
$write("%s",("\\\"\\\",2):f(\\\"\\\"}vtg=wxt;|bTaGV^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'3aqcC+bb.yZ6,*w-hbw-DtC+ftYa5?3rkiF,q=Sac3@|.x1uxof@E,KPRTEK2bjoVaR3i?v6C+A8kb?S\\\"\\\",2):f(\\\"\\\"{vNaSnbS/bhbCaDa4DXajuWalbj2\\\"\\\",2):f(\\\"\\\"{An\\\"\\\",2):f(\\\"\\\"{JoOtkQKLw7dKS\\\"\\\",2):f(\\\"\\\"}9b=4\\\"\\\",2):f(\\\"\\\"}A;A,*2bK=*Ua2kip;91sKYaxx@s73:Th?px=zc8@ipG|4|f>YYgIu<a,b*Pnp2:;Ge1aNNLTIv06yS2,7viwA6sKMr,bFZiBYv1hSKPv\\\"\\\",2):f(\\\"\\\"}Qcbz2f:\\\"\\\",2):f(\\\"\\\"}3a2b?r,9<6bbg7D,49Pc0?D?hbOadbIRw;01ltr=@WT/0x,btD<aME\\\"\\\",2):f(\\\"\\\"{b2|cBvx=F-bPsS4X-09ow5Dw20b@WRCYvfGDaP*6wc-\\\"\\\",2):f(\\\"\\\"{bhbOaX-k9qr\\\"\\\",2):f(\\\"\\\"{bdbL0Hv?EsvOjYvlo"));
$write("%s",("ZF:r5WGs13cmaprWaNa@\\\"\\\",2):f(\\\"\\\"{P|ybs3cOa.SjB>r;pdbRT1\\\"\\\",2):f(\\\"\\\"}lrXpB,e058@\\\"\\\",2):f(\\\"\\\"{U|clIh3v>qzUcbcA>K4vyZxEs9?aX-1+,KzWc?hbSCbEq>,b&6glb\\\"\\\",2):f(\\\"\\\"{sabD<oPM>\\\"\\\",2):f(\\\"\\\"}8Oa005bz30vW:BBEcPaFX?a1zJ,Fa-B*ZT/\\\"\\\",2):f(\\\"\\\"{bWaYa1bhbmLru6Y@LIUi9fbcbE-Pa.d<*yb:27bHW?aS-5b?afbzFawaRoEs/b7=t3Pu-BYaAa=y*qi3cuar?i-.bPa-P7C1bhbytTEr4cFbkb>U20SaDrNEujd<r?7vxKXn/b7qw8vt2bTuVvxK?afbkoBaGaT/7qQaUG6Y<y6YDZYa@axbA|ds+b?a3LGpEatf-AP*bbhbL4ybvb0v<zvq+|EKjS0v<z-;Pa2gI9d+bb+vCa-yZaJoS8kbGaT/8Fkt7=eZbzbevvf;sI|70T,Eo<acb3LGFvbuC7=1jNp++BaD?mbmCt\\\"\\\",2):f(\\\"\\\"}r\\\"\\\",2):f(\\\"\\\"}rFBa*bxbm;FX=akt-jK37+Ev78ir<ar3ldU*+v\\\"\\\",2):f(\\\"\\\"}vBf9|WC91<aUa.bPauCg:xqRSwbnpfGnWi-S\\\"\\\",2):f(\\\"\\\"{5b>i3s?am;1btLHq3Agf@av5zm*bItS\\\"\\\",2):f(\\\"\\\"}9rP864FaxbT94q?-i3crb=-@ay@dkl-TPI"));
$write("%s",("63lUaabkiJQ/>|b-r=QMQvuybLx.+ou/bPq+PQa=38/A0WaM\\\"\\\",2):f(\\\"\\\"{Ra/0/-hhHoZX1jMSV+dkNaZafgl|a|FfU*W12+M6Ux$6eIaUy3z:-T*<xW1jdIyw@FaZa.uB.rF*314wZ@Zfb/b?hbb0+6zOu-rv6C+jpC+9fxR=aUXsWagaxbA95/m3cycV3>r\\\"\\\",2):f(\\\"\\\"}2\\\"\\\",2):f(\\\"\\\"{rxbYaHE><>4p.==e9Lx-r\\\"\\\",2):f(\\\"\\\"{r=a,*W<ldo7M6Sa2hw<UaC<z+S1B-;KT*WCapfbStYPW4ey0b2bT;hbfP7bOC6b>wfPzbw=vbtuy<zbzb4bQaM6ysI9zqtBG5ub+Qgb**A?ogubiyCaCa5q8GqR4KJTG5ub5b>atbmb-VIzrz-rjp.4HquIkQJ7g:,7T*WaXq&6efbjbZpRNPaib1qQa38Ao.b,R||0bZqSuDImQ1qdysmS?R|*b9b?aSo-qYqkiWq-4A<dEXWQ<rztIC-PaapH4Ut+\\\"\\\",2):f(\\\"\\\"};^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^32^[2fha\\\"\\\",2):f(\\\"\\\"})3(f\\\"\\\",2):f(\\\"\\\"{#v3mja13(f\\\"\\\",2):f(\\\"\\\"{#,4353(|a3891(f\\\"\\\",2):f(\\\"\\\"{#(ntnirpn\\\"\\\",2):f(\\\"\\\"})4201(f\\\"\\\",2):f"));
$write("%s",("(\\\"\\\"{#)~4[~4bzc?iyo@JI*ISaAaySc<wbM/9w\\\"\\\",2):f(\\\"\\\"{@y@ArzbSaB;VaHEz@bbybYvfzxbYau@*InZR\\\"\\\",2):f(\\\"\\\"{tI0@Q\\\"\\\",2):f(\\\"\\\"{EaStV3tDK/Vaq<Waz|z@BYfzxbGa2Kc@QamQjb@a<xNaHEz@Y@ybYay@4N+\\\"\\\",2):f(\\\"\\\"}y.qzuwW>Vad<e<t;D-fGabk\\\"\\\",2):f(\\\"\\\"}?aVz+\\\"\\\",2):f(\\\"\\\"}K/n@yEVs4Nb1z+c-AGy,kiO==q\\\"\\\",2):f(\\\"\\\"}|DaOHa1=4+\\\"\\\",2):f(\\\"\\\"}K/:?Q8e2dCaVa-Iz@,9Rrxsn<P@D|Hw9-bSOaIRE|?aNt8*U@abqJW>60I62Bmq7w8b?aRU*wtbUaArcbiNPP+b<,T;=-@afbRuUG9O.bjdNa+bD,>SxhvN@aytpx?a1,@aIQ3UVzm\\\"\\\",2):f(\\\"\\\"}VaqCVzn|cb?|>SGaqAFa+/JhTrqqVzjb78Ya8g59ybDaiH<ajdeb,*2bWaGV/4JTmKPa6b|Fg21Zk\\\"\\\",2):f(\\\"\\\"{ybu?D+qxl2tsAocC3WZaCL55?u.U,bQa=aGtDIc,u=qINR4DPJzbDa@a/b9bhbAIujWaFXBaSazU3bf-I6PaVa><lbC<ebUtUadGg&b4<UtNa0D\\\"\\\",2):f(\\\"\\\"{b+b:T><7b=4z<u8AaOa@4Aa+bh@w<@a*b5b+y1b1uV68*TJ;0Qo\\\"\\\",2):f(\\\"\\\"}BFpDa"));
$write("%s",("=|Bat=TakinSZbK,AykbDaVap.Ankis4L+TuM4\\\"\\\",2):f(\\\"\\\"{x@B6wkq\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}cbSams~4azbTu=a.86I>aNunpy3KHNaxb+y1b*CebNHIo?fxHS4CakW3lNWPyhXKf5D.ZCv-;\\\"\\\",2):f(\\\"\\\"{/u|GkUXE\\\"\\\",2):f(\\\"\\\"}v+Aw7Cu=@g4bvby+tbL2zuQzW|jBbbYgpNSKTuGk<4c2aAaibu109Ot+>PXDMy0@u6R;xjNWaXp;qO-22@qbwUowxW.6h>bjc3+/b6RhyX,fx>a|LB*7CZ>38y6asU|r9R5mqdbcbn:1C\\\"\\\",2):f(\\\"\\\"}oXan\\\"\\\",2):f(\\\"\\\"{*Uu?NED|MpUaab>2Ra+e+b0q<=ybvb1|hEYZeEsvY3S0DiWadbcb,*Qald<F19?rd\\\"\\\",2):f(\\\"\\\"}S*qqebbbw|0by1hbRS:7a\\\"\\\",2):f(\\\"\\\"}lb<*O3aHbgb/q*4hb?aQyfbhtkd<FAwwyHV@Gx:0blbdK*qAo3qN+GP06\\\"\\\",2):f(\\\"\\\"{bOu*-PJ3E\\\"\\\",2):f(\\\"\\\"},kis4m77bPaki@o8D+b-Ic|-IQajA<aybZaFaRu0z?a@p\\\"\\\",2):f(\\\"\\\"{zO*?-dbcbnh-u6scbzZUarG,b>G6J1b296sUoKrfbxjmo2bYpE=eqaQa+b5D24\\\"\\\",2):f(\\\"\\\"}YZa5bG*M3aUb=ykqbb6scb=yvbkb1DTa1C58db6b"));
$write("%s",("3bBaD?sru?D+*3Q\\\"\\\",2):f(\\\"\\\"{*b6JqInJQ=SCdLbL+X+QQyFa<rE=\\\"\\\",2):f(\\\"\\\"}*z+EivbA:WabpvbwYKsKJ\\\"\\\",2):f(\\\"\\\"{z\\\"\\\",2):f(\\\"\\\"}Y5VPmtHOaKs*b;AWa\\\"\\\",2):f(\\\"\\\"{;2|XaVa.bk\\\"\\\",2):f(\\\"\\\"{0xf1\\\"\\\",2):f(\\\"\\\"{b6bPav3n@ibjmLrLOZa4AAoxxp59bT9Ao74>-HdrbV3=a=a\\\"\\\",2):f(\\\"\\\"{:nZy,ZaAoDs1Mkb+yFYP3|:F0ubm1bb\\\"\\\",2):f(\\\"\\\"}ZE=-b,bOtu4J|,bF4\\\"\\\",2):f(\\\"\\\"}bk9G5-tRNw<u=\\\"\\\",2):f(\\\"\\\"{:kb7bmterntmu@a7FF|?v6sXtRa+eDaq:66e|dp\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}JF;ttpJVWeHdbubr-6Jy,ub1bUx@aOo=6,R4\\\"\\\",2):f(\\\"\\\"}SC\\\"\\\",2):f(\\\"\\\"}DVa4@bbybj\\\"\\\",2):f(\\\"\\\"}<a8Fe\\\"\\\",2):f(\\\"\\\"{4b\\\"\\\",2):f(\\\"\\\"{Lu\\\"\\\",2):f(\\\"\\\"}4bx\\\"\\\",2):f(\\\"\\\"{xb4osXA.R|7+74lbvxufmo6@x\\\"\\\",2):f(\\\"\\\"{Aohb>atHk1CsU|nOox5H-;45Na:/bberSa|FScIoDaPXwJOwHLwbVv\\\"\\\",2):f(\\\"\\\"}JnM2CRnE|cBvq|tS0QEXzCoubG-3bS0Y00hCaW0p=Z:27r.U\\\"\\\","));
$write("%s",("2):f(\\\"\\\"}rr3babr.6qlbg2ab0hY0Va0yBa@aM;Owq3.bS0Bax?erSanMSaEo.dS0O<ixO<0bWsSaoPKMBam3W0p=Ctt;Dper(6e=aSaE=W:vqgIt<\\\"\\\",2):f(\\\"\\\"}qg|CoT|qM\\\"\\\",2):f(\\\"\\\"}Tf;E9f;R.7bE68CmK,b\\\"\\\",2):f(\\\"\\\"}bZ3kb\\\"\\\",2):f(\\\"\\\"}b4b|f/zc3imamKjbh6O\\\"\\\",2):f(\\\"\\\"{yb|be3a#cV?n\\\"\\\",2):f(\\\"\\\"{?7IwzAyb=a<a*bq;6:fbj=zt@a=pbIlT+d354bJA:siHb9<xXV57tHYv+dO/ts:E\\\"\\\",2):f(\\\"\\\"}|/rPa3CFaabC?tbz3YvYRpP:s3+sX4beoXwIoFCvb3C2VFar=51o=S*qSNpvbB,Rzk1\\\"\\\",2):f(\\\"\\\"}|0xcb>52-6S:s4bub5b7kh>8besubIMUasX*3Ao/b?N*o5HzZD=*o5DFzTaS,3WUawb,6e+d5bvbO/bb:8NRr|70qytsr|\\\"\\\",2):f(\\\"\\\"{C6b6YD=<-bb1bE6nxcAm\\\"\\\",2):f(\\\"\\\"{jS6t;sx8xHDZs>l|tbmb/*68W:<*<aR4x2UShbDaZRYaFYhb3UkqkiO=Z37b3bfP>akiN6?yU=QaSuqy9b*btqDA5sDa49\\\"\\\",2):f(\\\"\\\"}|c\\\"\\\",2):f(\\\"\\\"}+bOyFa0gkThO+@AaquC0EaY1FahEkbYg.;HOJt6@Oa-7mulbcbAwmxm;fgDz6xw|F"));
$write("%s",("a9>BaDKx\\\"\\\",2):f(\\\"\\\"{Ra80qAcbgB2vnZRS9r<7=1e>ZaXapT\\\"\\\",2):f(\\\"\\\"{1Fa9>kqc4Yi0.zbZb8bzb9blbiDRq=17C>xgWZ>3yzc<BWFYaGVu46f\\\"\\\",2):f(\\\"\\\"}dI>Yi70G-+Xxb7b\\\"\\\",2):f(\\\"\\\"{CXqZv2vhErNt3fS7bibvb\\\"\\\",2):f(\\\"\\\"{+vt2bM/VPQ<Raqux.3G4GHE?Tnh1htbG5S7ki5pt|NzB,Ta2h|f\\\"\\\",2):f(\\\"\\\"{ChbF\\\"\\\",2):f(\\\"\\\"{wbhbP|bbnKVP5bM4ytTqFi\\\"\\\",2):f(\\\"\\\"}r*b;s7u6Xd=>rdbMsAHrFUX5b,vc4o1.MhqZFvy=|0Sn5Au6b7vtb6b?aX:XFdbJLHL/bZn@s.r-7T*Itebn6n*hbDajb?u9s?aL9f|kbIrUo?Ls>ozUaCp498/rFFaWDfbgbh?6:OagfWz@3ZaS2L3<z0vffp\\\"\\\",2):f(\\\"\\\"}0b3boPXnPJub1*6fOaYanoXxOHgBf5E+gb8b\\\"\\\",2):f(\\\"\\\"}0fbGp>,kLOHhbAa7vh0\\\"\\\",2):f(\\\"\\\"}bD67bTqIw>2yZ9|mbiyeb+wzyUGzHnq;ivy+3ila6-M56YjbWat?3e>a\\\"\\\",2):f(\\\"\\\"}yZs\\\"\\\",2):f(\\\"\\\"}8bE\\\"\\\",2):f(\\\"\\\"}v+<xDar<=WC45?Wa1yur6qVr6YD<tbD6fyZ6lp+b<Lz+abq4i3aY2WaAoAJebzyFzzdCDfbhh9"));
$write("%s",("Q1NKs*wFa\\\"\\\",2):f(\\\"\\\"{qIA.b@IdbltEa9b\\\"\\\",2):f(\\\"\\\"{bcbo75b2\\\"\\\",2):f(\\\"\\\"{W|kbUS@JCY/3\\\"\\\",2):f(\\\"\\\"}|jsa|X,CwZY19jr>Ykb5?hbXuSwtjzbib-3jo\\\"\\\",2):f(\\\"\\\"{bzbiZ-Zjq2:J@=X?>>Vk+fb.8rgeb3+DKb+GaqUnwdbzbhbUilCVzFWmo/0tL>rjb-7@a:|8bJ4.86zZ*a,koYa.3S4<0ibNE**L|>o9|9xb\\\"\\\",2):f(\\\"\\\"}cb9s.4kolwv/jm9bNDc|0b,JykkbIw6YvbGP:t3Tgu.bfOebMue=5=?W8yfbh**ItbAaeCAz5OybgcIMYaqrmbkbEv5bzyNpabDKJARUzQN+h=\\\"\\\",2):f(\\\"\\\"{bJA<?Aw-3h=iIixcBV+CDPa@g2gy6WaMoCDS-Bs@smbBCQadW,bBaM66:cbwx@|5/VPNHkb+b38R@Nu6zL2Na.\\\"\\\",2):f(\\\"\\\"{A>FT?V6<s8DPnd?aCa*bEwxHo@6bFahrL54busabyba-7C/qsXPy:W/b;LWQVzSaSLEjSNdWlt1p+WN5WSGiTaRaDiS?cy8Ue|yIY<.vSa>a\\\"\\\",2):f(\\\"\\\"}boJb3YoOa-TStnqpupxlq:Wk.,t.btWlb.q\\\"\\\",2):f(\\\"\\\"}bYUlpTaGaU;qj|bUS1q,bbStq+AeU?ac\\\"\\\",2):f(\\\"\\\"}CaA\\\"\\\",2):f(\\\"\\\"}s>9w@3/Hv4;Agb-bsAzb|q"));
$write("%s",("abBa1b1,LrKHh?T*\\\"\\\",2):f(\\\"\\\"{x09n:2bkqM6S*IwmEl|ZVBH.bYO8bTaD6h\\\"\\\",2):f(\\\"\\\"}Ga<U8bbtHKc,\\\"\\\",2):f(\\\"\\\"}jjbH.|bjpnxT6M/4Bewaby0Oa|bz277Wi.b2:-1I@2:DTFa=zy4CDG9aB/xRacbrS64Za9s6qmbeb?aW>b,LxYUpr46|q:z?=ItYaorOSBfI9+oM/,bfbQ@.U5\\\"\\\",2):f(\\\"\\\"}lb5bWUkb58ApvGfqAq+bHqjSXw3U/Ois+JGaMqkSlhoIYadS4b:r-j7AnpAo1p>,2bquq,OyEvlb/bkimy/U7A7RAoubai:ro3tb747vYP0b1h38kiNIwb6L5KV6lb37s3EaU*2,jS2,Nq6=wsy3=|csTv|bPyTa1T9NK\\\"\\\",2):f(\\\"\\\"}xAq|,M>591z\\\"\\\",2):f(\\\"\\\"}AoSac<h<>7lhI9abiBTKdb>0477bjp4beb@l9<dM7<BRSCCB@4auVag2kiG,/|>aaSjbw=db<-2bbbuwPa\\\"\\\",2):f(\\\"\\\"}7Ccn:\\\"\\\",2):f(\\\"\\\"}w/yS<E-E9.*2gLxJSo5ubZqHs,SG>1jablb-tjS-b>akbYah?Nzd\\\"\\\",2):f(\\\"\\\"}AaNRF12h5gZ<lQrSKrtbG*wb70Oplby2L3UnL+|b6sUz@akQL7g:Btz3\\\"\\\",2):f(\\\"\\\"{bM5rS5g|uNa-bki;Q37FaG*>a|ubP>albtB<sPnQaY3<a1CAacujA>ttb09\\"));
$write("%s",("\"\\\",2):f(\\\"\\\"{bPa\\\"\\\",2):f(\\\"\\\"}k:sepYRvfZaSa0bSoAo6b7=SEXalbHqNE@Ckb:sxb>aPawktLSaP5CsJuwbJtPAUGyKfsNafb=aa27k4u.bPnv52:eMQB0:CP0voodsZa+b1RT|01243b/bSayHd<2bhbubYaWQc?Ovkb<04z2hBvpsXaMokxkbI1koA/M\\\"\\\",2):f(\\\"\\\"{*b3b,-HMUxRnyb8/q48b||A?tbW>gbA\\\"\\\",2):f(\\\"\\\"}UxfhMo3C:L8bs9=acye5qzpG:t4M8beb2/@G?a5bH>J/*Q\\\"\\\",2):f(\\\"\\\"}b9y|Fp?UxILJ1@3Io51kbJ/WsE8LxhOvz@L-dyyF\\\"\\\",2):f(\\\"\\\"{/l,@/|Q\\\"\\\",2):f(\\\"\\\"}J/fb6bfb1bc\\\"\\\",2):f(\\\"\\\"}Pa\\\"\\\",2):f(\\\"\\\"}owb21w<zu01U=izkbq0cbZEDa3bQa.8Wa,.g4jNjdp\\\"\\\",2):f(\\\"\\\"{@=i+1zGwbbAoabSa-b\\\"\\\",2):f(\\\"\\\"}bXay0L3vbws9bMrfPfbTa.*06F;kvf*VHONvbM6CLY;KOJ,\\\"\\\",2):f(\\\"\\\"}rfG/zt\\\"\\\",2):f(\\\"\\\"}=aEwQHf,;IYq9b2b3L9f3v\\\"\\\",2):f(\\\"\\\"}b9@8-8beg>q4oCaabnqisr3|.qGHh2u4bCacbTaY9\\\"\\\",2):f(\\\"\\\"{bQa+rkbIp3bkb1Cw?z\\\"\\\",2):f(\\\"\\\"}1bjD.5:pj9>p6p2<vryk?\\\"\\\","));
$write("%s",("2):f(\\\"\\\"}|:rrV3hET,9bbbrw5+|bCaapfw1u@yNpjbm5eg2qkdkhebN4Goub|-5bTak\\\"\\\",2):f(\\\"\\\"}u1C.7qN1.bJ1,|Rakt|Hs+/bnspq59Fp6bAovotoroSyS|ko<-?.eoh,boJ>44AaG5@\\\"\\\",2):f(\\\"\\\"{jb@yaKUvJrqxPaH2@<M6i5wt1-vbhcWJaMlby>k.S5Q5Hoxq|Kjmw@0ER\\\"\\\",2):f(\\\"\\\"}Rpaiyb\\\"\\\",2):f(\\\"\\\"}bj\\\"\\\",2):f(\\\"\\\"}=4jpgNtM5brMnz8bM;Ea2u49:Hj0mbC+j>4qa|,?O7ft@\\\"\\\",2):f(\\\"\\\"}Qr;Cx*|.1bC|jxK\\\"\\\",2):f(\\\"\\\"}.bDa\\\"\\\",2):f(\\\"\\\"{b@ItbHEO\\\"\\\",2):f(\\\"\\\"}abbb/b\\\"\\\",2):f(\\\"\\\"}wbbAaH2Y<7bD8FaIo@hAvTKUxOoMoGpUxEDOHjx1uf>5o+br;\\\"\\\",2):f(\\\"\\\"}b=aw?@aG7Aozb\\\"\\\",2):f(\\\"\\\"}bCa9+t5U\\\"\\\",2):f(\\\"\\\"}S\\\"\\\",2):f(\\\"\\\"}jF14ouAa71D?k|yy+bxjhj*b+-K;\\\"\\\",2):f(\\\"\\\"}bz+Fa4+PvlbiwMxgb\\\"\\\",2):f(\\\"\\\"}2tyowp\\\"\\\",2):f(\\\"\\\"}<zhD:io+bb5DYh-33,R:,3LkR\\\"\\\",2):f(\\\"\\\"{5?T\\\"\\\",2):f(\\\"\\\"{.1e61::lRDWJ@aQ\\\"\\\",2):f(\\\"\\\"}wtPaTox4t=EaRai-7o;qv"));
$write("%s",("uv6Ioab@=Qa<a8yp-hb.y7bUaM\\\"\\\",2):f(\\\"\\\"{/bAafxOj8bubOan\\\"\\\",2):f(\\\"\\\"{X|22,bF|1|2bjdJwi@s/mbn|Eao<9fL/2bEa*z1bVqbbJ6r9bbA4/bP5|FubS49b<J@ay>a\\\"\\\",2):f(\\\"\\\"}Ow/EOtP=N=0bL=Yg09RaKf+by,iB*bUa.\\\"\\\",2):f(\\\"\\\"},bf39uh6>K<KYvUt9D=aib*-Fa-bj|yK9bE|s?\\\"\\\",2):f(\\\"\\\"}b9bUa/bG=GFL@k1lwZaYakiK?AaUaeb-jLvibCa0514BaE7s\\\"\\\",2):f(\\\"\\\"{2b\\\"\\\",2):f(\\\"\\\"{bm|Q\\\"\\\",2):f(\\\"\\\"{2,7JNaUxIsYp8CEaFax;8g\\\"\\\",2):f(\\\"\\\"{oWavbQ\\\"\\\",2):f(\\\"\\\"{n|6blbCpTnYaH.WJIbTHI*nFlbdbT4:-kbs9YttD:sAo\\\"\\\",2):f(\\\"\\\"}j0b;qS2W;m?puo6+q-3=aiIGt8t=a@I1bQa*Iyb@a@aybfbFgGI1bfH\\\"\\\",2):f(\\\"\\\"{v=6QacB8hSaebyGeH|Gl2.bHqey+r7b5q.bFa>ao5tHZbY0E-5yaihtgr1bqGs1vtg:Ca>t?HS6o3*Icb\\\"\\\",2):f(\\\"\\\"}2R|>rm|6|>abk,Iz<Fa2*rg6bn/2Bgbebuq=a9bXa7oM5/l*bq0KHw+eb9bqs.b0w@\\\"\\\",2):f(\\\"\\\"{Xneb/\\\\\\\"\\\"),\\\\n(\\\\\\\"\\\"bWaSacbP?QaVa20VadyZa"));
$write("%s",("J|tbo49v/bW|i64bzo*bSa;qcqn.,b.b7bRaAGYaM5dyDaRauqu+kvCx-:d/MF*bsrki415b7bqi\\\"\\\",2):f(\\\"\\\"{bjb|bs,M,:wT*\\\"\\\",2):f(\\\"\\\"{r-ykiLsso2-9bOaIdEt\\\"\\\",2):f(\\\"\\\"{bTa?4kGJ|=|>a.bab<adbj0svqH5bF0?aS*azVzEaPa=aBaEajb\\\"\\\",2):f(\\\"\\\"}uvbY1y6<aGa6\\\"\\\",2):f(\\\"\\\"}1-EacsT,=3bbluME>azbybq;n4ebhr=DT?cAhstbHqKGG216K+RaebJ;Xa*bgkzbl\\\"\\\",2):f(\\\"\\\"}1>*b@|9b7bn/rxAowk5b/F|-q-NaZwsvwbq;\\\"\\\",2):f(\\\"\\\"}/t;Fa\\\"\\\",2):f(\\\"\\\"}jH\\\"\\\",2):f(\\\"\\\"{l,ixeb<a+b;p|E16lbfbFaqG46dtvbe0P-Ya*b|b,bVvQ8Na-,Va7+Fpq;a,yb-/PaID?|zb>aO*DawbL\\\"\\\",2):f(\\\"\\\"{h-ib\\\"\\\",2):f(\\\"\\\"{b.3Ss1z*t8lKFvpPD:xAa=azbdr0vTo.3+v,-pzz\\\"\\\",2):f(\\\"\\\"}nqUadbb3j|?C?aFa6r1Cft|f+b<==DZa1CibybOhx/Yhcb:+F|z+<t=69o2*o|.hbbi\\\"\\\",2):f(\\\"\\\"}FaNCibooU\\\"\\\",2):f(\\\"\\\"}H:pDMumbZE7bCDQag-<@N>Saf-\\\"\\\",2):f(\\\"\\\"}qV>xs/b\\\"\\\",2):f(\\\"\\\"{bNa<xwbguTac"));
$write("%s",("bmb/@-7?|q,Oa7u5uFabqKoY@hb>o8bqCSkXao=tbTqBa71R\\\"\\\",2):f(\\\"\\\"}Y?*@\\\"\\\",2):f(\\\"\\\"}+Es/4Ua7b>?Ez7\\\"\\\",2):f(\\\"\\\"}ZDCp8g4bD,xbEaUa:pR>vzR4XpirYahbAoh7YaY310KCO@ibY;:05b2bAo6xOx8C6C,uWax8.1.:,\\\"\\\",2):f(\\\"\\\"{OB@lMBwbgbl?Yahx/y49/<1u/uh,5bdb846p85*\\\"\\\",2):f(\\\"\\\"}hb2b6@8DKfebQa88ZoUa?a8bIs=amb,*tbNtR|<9O/jbmb3|GtzA3C8A-u.43b7z5zr\\\"\\\",2):f(\\\"\\\"{F:5b?<|,O*Z3/bvbwbD,*by,r9Daw5G5Vrr4|bvbubv8BfkiB1isOhOa5720e3l,L@q,h@@a4b1*ib/b5bSa|b<a-vzdVpM+V3ibabYa,zykbq3bVv4brwp\\\"\\\",2):f(\\\"\\\"}2|S<i2/82*R3Us\\\"\\\",2):f(\\\"\\\"}b.xVz/b9+kdNaytS@iujpS*8*yb;pPaUa7sctub-bdlXBF\\\"\\\",2):f(\\\"\\\"{p16b@2t\\\"\\\",2):f(\\\"\\\"{Xy+bI>p+:2Csvn2:r8d*G@=lE@6b*=xbZau1T,rgf+N3u\\\"\\\",2):f(\\\"\\\"}/4:/59+bNaVz*bRp|bpzBaZsSnN+OaluZaKf=oJAixWaP*fhy<ibzbkb:q2*Va|3Y0+x3bo<1bSzNkI,g;iwOyubFa\\\"\\\",2):f(\\\"\\\"{b+vYabq**Ht/b-7"));
$write("%s",("\\\"\\\",2):f(\\\"\\\"{bTrtlq7D?\\\"\\\",2):f(\\\"\\\"}+MA7=X,?a4pzb1bPywbP*N<-bfbr=3qp=Q10bNaS*;AdY2oG*jbL=3b>a+|h7\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}2b1b<,f3yb-jv|u\\\"\\\",2):f(\\\"\\\"}1bl>DrS=bb3+e9Aa0bbbM>S2hbps8z+bbbki<1Kzo245rr=;y6AaL0e00r-buyzb+bXarzAuhb7=1bisjb,b6b-bWaAaebCaL<,b.1*1@>@l>>2:<>q,VaGw*wp\\\"\\\",2):f(\\\"\\\"}ybAavbOtEor<@aZaViDa+\\\"\\\",2):f(\\\"\\\"}WaAq3bG\\\"\\\",2):f(\\\"\\\"}mbbb46-;ubXambGiez1hwb@aebcbJ,<x9sczD?inVa?aWaV?4uzqqu@aVaNhAoWaqzk.?a9?cyJ1z<4bkbU0>aAox7g.Vav8+yWaV38b=5>ayktbp=J15bVabbgbgc,babPvjbj43bQy?.65457bec\\\"\\\",2):f(\\\"\\\"}w-bwbdbAqu?\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}J-49|?lt3zY\\\"\\\",2):f(\\\"\\\"{@uM,Yafb\\\"\\\",2):f(\\\"\\\"}b3bu*BaQaN1EaG5|,-b?avtsmOaxbybA=Oy598bS8DaabQ16xXatbSs5\\\"\\\",2):f(\\\"\\\"}==i9iw1up/2uAad,y>FpUa>plb49,qXp,bkvf/8<=lb*.15<N-jdlb@\\\"\\\",2):f(\\\"\\\"{ub>aQamzr3|4R"));
$write("%s",("ae|/bLpJ:guj4hbIdq=@9d3hb.b\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}a3B*E\\\"\\\",2):f(\\\"\\\"}Pas:Ho5/Ho0bO0z9T,;rU6vbb;eb-y*bXaAoDaAwsmKrWas/9bPz,bGzNt6p\\\"\\\",2):f(\\\"\\\"}b8bm\\\"\\\",2):f(\\\"\\\"}RaZa3b1uko*o\\\"\\\",2):f(\\\"\\\"{ybb|b16;ptbjbAam7Tafb@xhy=aOqAowbbwkt+0x9Kw,*2hi,TaSr/ykb3yMoy1>axb>oyb0bOaPa5b.bcbxb\\\"\\\",2):f(\\\"\\\"{b0b2<0bT,kb25jpQa?a;x|bk9Np;y-bmbTvFa3y,-OpTa>uzcsw+b@aD,mb=4Uv1<t;h<Uav8WaEaSak.PnWaWaB-D-xo=lb/d6.1/:o8Aam8Y9Ao1wz+\\\"\\\",2):f(\\\"\\\"}*h<prr.TyorTa=aWakbfpjbvqK-ibDa2gVaHpWaTa@aiyvqe<s.TaBambB-PaWa=4EaqyCaibn:kiM3wbGwvb=oPs3bw+lbAw=95b8bxu@-ubdto*Ya4bUiv|N7lbKwnuw4/z\\\"\\\",2):f(\\\"\\\"};=6<6ZoUxUye89-g2Ptkx-v5bjd>ac4fgwbzb6zwk?a0bZoP*7bl\\\"\\\",2):f(\\\"\\\"{<aAocbN7YtYaNkW0.l3bg|0b,bF\\\"\\\",2):f(\\\"\\\"}mb3zOtOalbyy7bzb>yXafzquvu/b\\\"\\\",2):f(\\\"\\\"{+|b?aNuLp/booT\\\"\\\",2):f(\\\"\\\"}R\\\"\\\","));
$write("%s",("2):f(\\\"\\\"}9yfg9r9-Sop\\\"\\\",2):f(\\\"\\\"},b=aY8-bW8P\\\"\\\",2):f(\\\"\\\"}Naj-J9kbczPalb.1C3c/F3c6D3ovq8|1*\\\"\\\",2):f(\\\"\\\"}y|z6>ajbUi3rBav:ib75\\\"\\\",2):f(\\\"\\\"}bL,J6Saix|4Xanpvbgs<9a2z2FaAoVta,*bexFa0bvbgp1\\\"\\\",2):f(\\\"\\\"{j+d3jbpjhbrgj7+oXa**Xa\\\"\\\",2):f(\\\"\\\"}*Gg|b4tab2tVaZu:|hbPa3bB\\\"\\\",2):f(\\\"\\\"}@\\\"\\\",2):f(\\\"\\\"}=ayb/bfbw8Z-PnJ8tbTaww7blb>aJ|@aW5Pa0vybSaFjI\\\"\\\",2):f(\\\"\\\"{G+OatbJy.rJ8=a1bUa8|BaO\\\"\\\",2):f(\\\"\\\"}F|\\\"\\\",2):f(\\\"\\\"}/V8TaDaEaAoUoA*ubd.Nufb1w/b\\\"\\\",2):f(\\\"\\\"}bj045hb8b*blbPu?am3Va6zjb+8/hkbj0jbIq/8lbyb@y3gOaJpo44bSa\\\"\\\",2):f(\\\"\\\"{b=oCaXa1bjb+bjb,*Dao4Gi:.zbNaXy<|jb>7DaJ1Ar1bSaPamblbVakvG3-\\\"\\\",2):f(\\\"\\\"{E38,a6VaOajxYaHpp\\\"\\\",2):f(\\\"\\\"}Aoa|I6v|/bEa@a+uO5t\\\"\\\",2):f(\\\"\\\"{lb+/8yS*:tOa<ar\\\"\\\",2):f(\\\"\\\"{*|Pa?a;7Da978bwxjm\\\"\\\",2):f(\\\"\\\"{b+o+bUuc2<7zycxOa,b<aRay6xh2bkx46K"));
$write("%s",("tFaa0RaIo>p;pw|oy7b7bebL0lbjbruG5dvhb,b\\\"\\\",2):f(\\\"\\\"}rBaF|ibvzQaw|Xamjibt-r\\\"\\\",2):f(\\\"\\\"}PaJ.0bubU+Lqy6Q614Tq4bbwK6I6Fa1b<aVzW16z3*bxvbzb46QambabmjSavbgb0bFi\\\"\\\",2):f(\\\"\\\"}bxbIp=a3zcbgbzwzy2b<aiucy>aFaBfCuvbRaBa-yczF\\\"\\\",2):f(\\\"\\\"}e3L\\\"\\\",2):f(\\\"\\\"{Gvq6Ratbwb\\\"\\\",2):f(\\\"\\\"{x3zWaCuzo.b\\\"\\\",2):f(\\\"\\\"}b5g<avbQaNa7g4bltVa|b:+.\\\"\\\",2):f(\\\"\\\"{:,Fx.\\\"\\\",2):f(\\\"\\\"{DxB3\\\"\\\",2):f(\\\"\\\"{0r1@5Za>5lb*odbXaGp7byb.b,bAaub?ofbF\\\"\\\",2):f(\\\"\\\"}kb\\\"\\\",2):f(\\\"\\\"{/@z:+mw/-f+/y35Aak.9bub0bQ\\\"\\\",2):f(\\\"\\\"}bbxbqy6bZalbquVaAoq|2uRp+o=rbp9rQoL*Dp,*EaybxbAflbxbTa24kb,b>aTahbLwX|cqubG.8bdb,bf-y1m3cbMyE04bKz2b/bUa1b?zxb8uIo3bbbmbjrVs3bLo4b\\\"\\\",2):f(\\\"\\\"{dIpDaT0mzRaVa\\\"\\\",2):f(\\\"\\\"{vSa0p4tl\\\"\\\",2):f(\\\"\\\"}r3Qa8bjb<agbBv,b8b,okb8b8bUzhjyb3,Oak3xbXa/blb6b2bytQaTaCadyFa<aabgugb=a8bx\\\"\\\","));
$write("%s",("2):f(\\\"\\\"{wb\\\"\\\",2):f(\\\"\\\"}b\\\"\\\",2):f(\\\"\\\"}0UoPak3A2kb\\\"\\\",2):f(\\\"\\\"{bfpX-AoCaWa\\\"\\\",2):f(\\\"\\\"}b*bn|2btjAo3bZadb\\\"\\\",2):f(\\\"\\\"{xdbvn.1e*Ex+1/\\\"\\\",2):f(\\\"\\\"{,10bmbvvqo|bN\\\"\\\",2):f(\\\"\\\"{ebzu,bGau\\\"\\\",2):f(\\\"\\\"{foJstb<al3zwNaubcbzb/bBafbkx1bu1lb.blb.u0bTz+bkbQa9b6bDaebzbj\\\"\\\",2):f(\\\"\\\"}fbTuWaVqZaBaxbvb7bDacb>0bx=roz>aVaBadb3bk|.oqybqlqbbj0bbt|xbbbTaX+Vp02.2bcQaohNaNa|b@akb<a|ba16bmqosz|Eav+ib1bj-fclyjbIv-b\\\"\\\",2):f(\\\"\\\"{vGaRxDa5bcbi+U*w|@aFaYaArPaZp8bcbVa=aUa<p3bM,K,6z-broZa<albt,Rakq6z9w7bv*Pafpb0\\\"\\\",2):f(\\\"\\\"}bGur\\\"\\\",2):f(\\\"\\\"{F1gbjs2v?.kblw?1=1\\\"\\\",2):f(\\\"\\\"{b2j>aMsAaAoOaa\\\"\\\",2):f(\\\"\\\"}Ohdb21TanwAofbq-2b.qwb4aY\\\"\\\",2):f(\\\"\\\"}Z\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}1a*7,e/mbjbPa.bY-3uJ,yb5r1b+b>o0b6\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"}oubt\\\"\\\",2):f(\\\"\\\"{wbRqOtzr5bAaPa*"));
$write("%s",("btuPa8b10eb7|Ba<0vbUafbR-U\\\"\\\",2):f(\\\"\\\"{Mhmb,|Tp3beb>\\\"\\\",2):f(\\\"\\\"}AahbltfbXadbbb\\\"\\\",2):f(\\\"\\\"{b,bXahxib-iwbVazbG*Gaeu+bBvzbfgAaBa+b*b7q<,Zakqdz?aTaVnv|4binCsdbfxX,;xh,Aa7xibm\\\"\\\",2):f(\\\"\\\"}*bLxFg7bjdibebQy\\\"\\\",2):f(\\\"\\\"{bfbEadb\\\"\\\",2):f(\\\"\\\"{bL,4qfbw+MvkiN/?ykii|mbAo|b2bjbgbgbzbC/9bfqWn1,Ca|/=aNagbRaa-B,+bRagb.bhy0q>a,tNaabE\\\"\\\",2):f(\\\"\\\"}F\\\"\\\",2):f(\\\"\\\"}s/i.?aX,gb?|@a7bBa3bS.fbW.CaKtD,>a7bzv\\\"\\\",2):f(\\\"\\\"{bDalbGsOar.>a<x7bvn\\\"\\\",2):f(\\\"\\\"{ia/tn6,Hx9,6.4.RalbZ,3b=aSa=a/bb.QaD.a-G\\\"\\\",2):f(\\\"\\\"}=aabG\\\"\\\",2):f(\\\"\\\"}4bzb8*Kyk.6b0bjbrz=aUt?a+bebZaD-wbhp3bibizDar.<aWab.lylbQa/hVap-RaD-OyVaPa>aEaAaZ+1hRaWaUaVy=aEalbgbbmb.TaSa@agbNaL+Ra.bSadbxb.oE|t-0hYa0v=agbUaEaB\\\"\\\",2):f(\\\"\\\"{mb@aRagpUtCaSa.bRa@aWaUt6bjb.bYalbabXaZa.bF\\\"\\\",2):f(\\\"\\\"}Na<ths4*FadbVn1bL\\\"\\\","));
$write("%s",("2):f(\\\"\\\"{j\\\"\\\",2):f(\\\"\\\"}db9x0b1qOaLp1bibUa\\\"\\\",2):f(\\\"\\\"}b?aJySaBqxbRa6b,ts+Na@aQa6b*bboBa\\\"\\\",2):f(\\\"\\\"{bbbjuOa.bCa?awbabFgLxv\\\"\\\",2):f(\\\"\\\"}Bajbzb:thwAaykmbBawbUagbOx7v2bVaUaR*6bebR*ly\\\"\\\",2):f(\\\"\\\"{bZ*?akv>l5,\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{rnc*X\\\"\\\",2):f(\\\"\\\"}PazbRa-bR*T*SrbkRojb0bVa9bBaVaFaRa;yN+L+Py7+xq8bs\\\"\\\",2):f(\\\"\\\"{@a;\\\"\\\",2):f(\\\"\\\"{DiOaWa.b*b7bXqZa>a-bXa?aOa=a3|0b?aeb8b-w7rcb8w3+cbwbSalbPaldIvkxhsauEaXaOaykepwtUtykybCa6bXaUahbjbt\\\"\\\",2):f(\\\"\\\"}Ua4bYaDaubWaxjqueb6bwbF*Pa1wmbgb\\\"\\\",2):f(\\\"\\\"}b<wcb\\\"\\\",2):f(\\\"\\\"{b=axb6bVrTr3bDaUa\\\"\\\",2):f(\\\"\\\"}q*bjbOa3blyCsVa+b1bVsUaX*Zamszb4y=oZakbNazbYyPa1bwqSrib7oDrBaslAa,b\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}DaUo\\\"\\\",2):f(\\\"\\\"}bab+ohs?afwbbCaki5*Ra+bAo0bib5bZaTaPatblbOa0bOw|bRaxbtb\\\"\\\",2):f(\\\"\\\"}beqxbx\\\"\\\",2):f(\\\"\\\""));
$write("%s",("{tbrxcbYa<adtEa8bkbBa4b\\\"\\\",2):f(\\\"\\\"}wBv\\\"\\\",2):f(\\\"\\\"{o<avn.\\\"\\\",2):f(\\\"\\\"{/sonGx*\\\"\\\",2):f(\\\"\\\"{.\\\"\\\",2):f(\\\"\\\"{|\\\"\\\",2):f(\\\"\\\"{+\\\"\\\",2):f(\\\"\\\"{z\\\"\\\",2):f(\\\"\\\"{ubzbwb7btbebhbBazb+v8bbbkbXampE\\\"\\\",2):f(\\\"\\\"}Raab1bt\\\"\\\",2):f(\\\"\\\"{luq|QavbabcbKwr\\\"\\\",2):f(\\\"\\\"}R|>wh|<rkiG|gbjb9bvb5b*wDa=tot5u4bfbOa8z6uOasw;w9wOaTaub9bxb?xcbhb0bdb-bOaCazbubkb*t\\\"\\\",2):f(\\\"\\\"}|2bYaNa\\\"\\\",2):f(\\\"\\\"{bZbXaXaPaKxYa|bmovbfoFa8bro8|cbkq*bGyAoFaOambmb*b+b,bOa/bjbjb\\\"\\\",2):f(\\\"\\\"}bNrubZaibSaj|7gBaUaYaQa3y*b+|\\\"\\\",2):f(\\\"\\\"}|eb\\\"\\\",2):f(\\\"\\\"{bgb*bibRsOa@aW\\\"\\\",2):f(\\\"\\\"{tbabfbwbmb/bybruogVa\\\"\\\",2):f(\\\"\\\"}bSaubAohcXaTavbvbXn|b>2iytb*bAafbebsw4b?aUa8bvb0qdb1bcbvb\\\"\\\",2):f(\\\"\\\"{ryb*bmb@ukbsrywSaWa;p=ahy2v5rUatbxr+bUv<atbSavsxsvszbkvlv\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"{jv.sIx,skv1s-sBx2jNat\\"));
$write("%s",("\"\\\",2):f(\\\"\\\"{NqPo@aab8bfbbbqs4blbXa>aWzUz+dYz6qNabb?qjbJvZqabRaUaNadb2bPa-bdbTa+ukbebxbWaIw9b9bab|b7bxb\\\"\\\",2):f(\\\"\\\"}qvb-b5bRscv-b/babQa/ubb.rOahbabtbQajb\\\"\\\",2):f(\\\"\\\"{b4bhbCpxbAa.bpy0bAaab-voo;iCasswb5y8bEaub\\\"\\\",2):f(\\\"\\\"}b|bWa4t@yRafbQaAvVa8bwbkb6sAa2vUaOaIymbfwebSaiyPawb/b4bZa=aOa>a?aKrzb*o<xAolbapit*bhbcbEa5bYaxu+b>assOwRakb2bAufb3bTaabibVaYaVa<a6btbgb3b,qabTa3bfx;v/bDa0bfbOxdbUavuhjubdbIqXafb8b\\\"\\\",2):f(\\\"\\\"{bBa8bEwAa1b|bpxgb9x<oNxYw+qAo-bAatbzb\\\"\\\",2):f(\\\"\\\"{i\\\"\\\",2):f(\\\"\\\"{p|pyizpkvmvkvnvibEa0b\\\"\\\",2):f(\\\"\\\"}b9xCaxbib3bKs\\\"\\\",2):f(\\\"\\\"}bmbUaDvDaytZs-bOtVajpwbebbp:tvx\\\"\\\",2):f(\\\"\\\"}b=opx7b>aNalbvjgb|bPaub*o=a*bru/bXaeb-bStab9b5b1bAo+b6bTw6bPrGt,b:rwsNaOayrXahbtb7b0b8bmb1b-b*bOa-vlbib>avbebPa4e*b=aYaRa9bTatbruWsgbTaAaWaybAixj\\\"\\\",2):f(\\\"\\\"}b/bZa*"));
$write("%s",("bvo;s4b,b\\\"\\\",2):f(\\\"\\\"{bXa9rRaUi=abb@a0b+bTagbwbSuubabZabmTaxbkqdrBa,bZskbArsvQa0b=a5qrm;p5bNarv\\\"\\\",2):f(\\\"\\\"}otbxj,bZa6b.b*q\\\"\\\",2):f(\\\"\\\"}b\\\"\\\",2):f(\\\"\\\"}bTaYatb5vcb-tJqkoSaKsEa?aAoZo/bdb7bZa0bXaNtYabb6b\\\"\\\",2):f(\\\"\\\"{b1bdbAa@a\\\"\\\",2):f(\\\"\\\"}bAowtutNaKfHqXaqr/rkv*siv+s4a0s<l|sfbRnBagbxbmb<a*oPaCa.bAivu|bDa1bXa/lxbeb5bEa5r3rRs*bEaCayb8bhhRaBftbdbYa3b6q0gWaooPaXa6bibmbxbgbkbab*b4b*bwbFaUaUnFacb1b7bxj8bKoDa2bmbTq8bWa0b9bmb0bkbXtTa\\\"\\\",2):f(\\\"\\\"{bOt7bkiBr2gAo@ambEjSaSaXiVaSa3bYa:p=tab\\\"\\\",2):f(\\\"\\\"}b+b/l@aAa3bPa|b6bht?a/b-bRaqswb>pEa1bWa8b7b4bFgEiRaujXaHoAfYrdb=q7bNa.bCsxbCa/boh-bAombwb1b2pdb+buoUsvb\\\"\\\",2):f(\\\"\\\"}bzbTaFa7bSakbFagpwb,d6b>a,b-b\\\"\\\",2):f(\\\"\\\"{bubfbzb@aXa4r2rQaXa+bGiibAoYaeb=r4bPaxbFa/bPa+bfb+bFa5m\\\"\\\",2):f(\\\"\\\"}ryo1bfbSa8bvq.bmbhbQaprvnyixp"));
$write("%s",("\\\"\\\",2):f(\\\"\\\"}syp\\\"\\\",2):f(\\\"\\\"}pwpvnvnMiqpUaVa5bRaXa.bZafbibfqbbbbQaUaAaHpzbWaXabb3bAabbcb\\\"\\\",2):f(\\\"\\\"}b@acb1hvbjrUa,bTaNa5b3b,bAoyoYaFa|bmbRaub<aVaIo5b@aAoebyb3hvb.bib6bdb5b/bZq7b3h>a8b.bTaYq=a6bkb-b8b2bFaebOaYa0bwbyb5bkb5bOaubQa\\\"\\\",2):f(\\\"\\\"{b.bUaSa<aubjbcb9bzbjbRazb2b@aSojdQalbAoVa>aXacb7bfb-b3bUaki:oVa0b/b7b2b*q|qzq*b6b|bUavb@aublbvbVa\\\"\\\",2):f(\\\"\\\"{bbqib,bdbFa\\\"\\\",2):f(\\\"\\\"}bkbdbgb4bTa+b7bdb0bPa,b7bwbAo,blbUaQa>aibSoTajbTa/b0bWaBaFa+bEawb6bSaXa\\\"\\\",2):f(\\\"\\\"{bebmb+bDaFa5btccb0pFaDazbEaEakbbbfbZajb-bEaabjbhblbYaZaqoDaDa\\\"\\\",2):f(\\\"\\\"}bwbQakbcbibvk\\\"\\\",2):f(\\\"\\\"}b7gAoNa,b2b|bhbNaBanpLhhbwb\\\"\\\",2):f(\\\"\\\"{isptp8lrp8lupun\\\"\\\",2):f(\\\"\\\"{iynzn\\\"\\\",2):f(\\\"\\\"{ixnvndbDakbRaCa0bZaCa>aOa4bUazbCaebwb\\\"\\\",2):f(\\\"\\\"{bybib+dcbbb,bebYaAo4bDaYadbebXaBaabwb*bCa5b|"));
$write("%s",("blbGa;ogbvbNa1bkiqb7b<a>adbCalb,bYa.o/o-o+o7b/bYagbibjbDavbDaQaEa+d0bybeb.b-beblbzb,bNa7bvbCaEahb<aCabb*b8hQaub*bWaQagbSa,bEa7b6bAaEaXlBn1nJm\\\"\\\",2):f(\\\"\\\"{mym*nXfMm-m<n;afn.m?a,mfnLmJl6n-bXlCmCaIlcnwbicfnKlxm-nEaimMmzmIl3mumsmvn@l@lpn4asn9ayiqn8lnn;l\\\"\\\",2):f(\\\"\\\"{i?l/b\\\"\\\",2):f(\\\"\\\"{f-a;hub@h8aDmQm4mVmHl9aEaOaMmKm<m2i:a-bMm=aAa-a=m7mCaimmm2m@a<a-b|e@m6mamwmlmcmamYl*m5m:aCa|e/m>aAaxmhmcm9aFldmAa:kTl|evm/lXlkmBa-aZlSlQl*bvbtb/b-a+bIdLlemMlVl@aTlXlSe|eRlWl?aAaIl\\\"\\\",2):f(\\\"\\\"{bGlNlLlFaJlHlFlHaDl9a|eElxb8a+e-a1beg8aXf,l8arb|eidxi=l=l9l3aLiyi7l-fziylOhFf6b-a+czbxbubHaqb6aqbEiFiDi5aqb@g-a,bAfzb.bKfnbxb\\\"\\\",2):f(\\\"\\\"}ikiZgXg\\\"\\\",2):f(\\\"\\\"{gag\\\"\\\",2):f(\\\"\\\"}h6hjk7jqk?a=aLi;dLfbk7i?kvh=ktcBa3aPhIgDiwbPf?a@krkWjBa?aKi6e;hrbck7hDhZj*hXjDa?a>aKi2b3bGiUfyj8f2i-bCjCa"));
$write("%s",("3aKa\\\"\\\",2):f(\\\"\\\"{b;a3gwbccIa3b1b-j,b|b0avhakik5jCaKi.bti7hvhQiOiMi@aKiyb3bTj?a9j5i5h6jBaLiMf1i\\\"\\\",2):f(\\\"\\\"{g\\\"\\\",2):f(\\\"\\\"{gsbubwbki-aDjBj:a;b?j1b0b-b3aAa3a7b-aki.a:b:b,b7hWhPimiNi@a3a;hwb+b-aPcuj/b8b1bPcxb;aUf-b:fZapg|b.b5b-amj>i3bWfvb|bIgGipgfg3bgf;a<b:b3b-a8bIg,bxb2b2btb;a7h*h6iPa4i3a>a3a5anb-aEi/b3b4b.bHa8byb2b2gtbWfxb5b+bYg7h5hliYhWh;d+cKfHa-i-iFaGaji|fld4a.gwi/auh4a-afgdgMaFa=aWh-bYhDhChGa+bJdRh9a/b5a|fCc8g-bPaBaobDhHfMa9aMaIa5axb3b.b4b0bxbzb-btbeg7hkg5hGaMbHg2bzb;azbLfccJa7b?a?auh*hCdYaOaVafbVaibNa=avhvh?a;aSgVaNaUa.guhkgvbpbEa*c7bEaBa>aDa>anbJdubSczbPfIcQgyfwfuf2bsfNd3bHa?e-a-fZf:aIa+c9f:avbldub4bcb-b3ggc0gHaebdbJaGagfef8a1bxbwbtbxbUaac|b3bdgfb/akgzgtbxcRf?a1akg-a6a5bhg>azd:a,cNahgwb.b;b>aagob,c:a-a.b\\\"\\\",2):f(\\\"\\\"{bvbxb5a1aob,fCe2b-a:b1dtbHa6"));
$write("%s",("a/c2b/a,fPcFf/b:b6aKa6e1b4eIa8btb1b1bNaGatb5a+ctb,b-a\\\"\\\",2):f(\\\"\\\"{fyb3dMd-aDdBd@dmf/aob5a.d,d*d-b4b7eSc;axb+b.bbcZb0cbfJasdHa/aed+e0cGb/d,btb-b4aWbudpcgdLc=chchd6areOapc0cNb/a;bje/eGaHb5dedOb.a8aNd8aLdLa=a>aIa\\\\\\\"\\\"),\\\\n(\\\\\\\"\\\"OaJapb6a+e5azb+cdcfbhc;aOaFdYd6aHaCa@aIaQd8aHa=a.cIbCbMd\\\"\\\",2):f(\\\"\\\"{cycvcocRapcXbocTa;b;bpbgbYdJaGbRanbQaJagbnbcb>dqc5dpbebnbOa8a0c4aJaTa5a+btb5bxbJaQa,c*cRa5a1bzc6aedMa0c3bldjd;aeded8ard5a6a5aedxb/btbvb2bxb,c1b4b3bxb1b0cocPa8aNapcMagdUc3b|b+b/b2b4arcFbnc4a=a?axbtc4aSbJcPbKckcic+bZb3b-bzcXbqcFb5aMa/ancvc+b+b|byb4a9cVbNa5aRb7cFbnbFbMapb2c.aMaFb.a4a5aJaOa-a-b|b-aeb5aicybHa<b/akc>a>aXb6aOb/a8a6a/apb4a1b.b3bvb4b1b3b2b-b.bvb4anb/aJaPa5a8a4a6apbEb5a5aBb,b9a4apbpbnb8anb4aGa=a:bJacb!\\\"\\\",2):f(\\\"\\\"})46(f\\\"\\\",2):f(\\\"\\\"{#~[2xha=s,y=z,13&X"));
$write("%s",("3^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'yay,]99999[gnirtS wen=][c n3aea\\\"\\\",2):f(\\\"\\\"{)v]y3b&a(niam diov citats cilbup\\\"\\\",2):f(\\\"\\\"{RQ ssalcz4rfa cdlnl3c/a;maertStnirP/oi/avajL tuo/metsyS/gnal/avajm4bdateg@3doa2 kcats timil.v3dga]; V);Q4aC3ecaL[b5aX4hha dohtem?3e;4nga repus&3ecaRQ@3cgassalc.<5joa(=:s;0=:c=:i;)|4ajaerudecorp/3fqa(tnirp.biL.oken\\\"\\\",2):f(\\\"\\\"{.3bianoitcnufR6\\\"\\\",2):f(\\\"\\\"{sa(rtStup=niam^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f"));
$write("%s",("(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^32^[2fha\\\"\\\",2):f(\\\"\\\"})3(f\\\"\\\",2):f(\\\"\\\"{#v3mja13(f\\\"\\\",2):f(\\\"\\\"{#,4353(ga36(f\\\"\\\",2):f(\\\"\\\"{#j4[j4boa(etirw.z;)tuo.N8aba(67b~auptuOPIZG.piz.litu.avaj wen=zG4Zka91361(f\\\"\\\",2):f(\\\"\\\"{#tm4[m4c5aR0Z0Z/512152353/2/2166263=4/3141726??:1518191:1/@4[@4cda*6 Q5[p4dea1312^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'5[w8[$5ofa41310r4[r4c7=[B>[j4[^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\""));
$write("%s",("\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'6pma(amirpmi oicy4[(5[j4hma++]371[]591[?6[?6cpani;RQ omtirogla\\\"\\\",2):f(\\\"\\\"{4[\\\"\\\",2):f(\\\"\\\"{4cua;t:\\\"\\\",2):f(\\\"\\\"}%%%%\\\"\\\",2):f(\\\"\\\"}fi\\\"\\\",2):f(\\\"\\\"}*-84\\\"\\\",2):f(\\\"\\\"})48z3b(a]i[\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"}+17\\\"\\\",2):f(\\\"\\\"{<84.;i:-i602\\\"\\\",2):f(\\\"\\\"{;i:911\\\"\\\",2):f(\\\"\\\"{;j:632N4Zsa7218(f\\\"\\\",2):f(\\\"\\\"{#(tnirP.tmfIIcfacnuf;&4[&4bdatmfn4[n4cgaropmi;ILagagakcap~4Zea1304T6dbapD6[r4cba-l4[l4bjatnirp tesY>[ca89&AafantnirK7[ia959(f\\\"\\\",2):f(\\\"\\\"{#fp4[ga^64^\\\"\\\",2):f(\\\"\\\"})74[8awa,s(llAetirW;)(resUtxeT:Paca=:R6[ba1Q6ak8ap4[p4adaS Cn4[vEaca&(z5[z5aba 06[06[06piaRQ margo^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\""));
$write("%s",("\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'5[t4cjaS D : ; R-5[%L[j4[j4o%6[k4aqa. EPYT B C : ; Az4[56[j4[j4nka)*,*(ETIRW/6[J7chaA B : ;s4[s4aba [2cr4[*5dia: ^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"' ohce4B[ka3(f\\\"\\\",2):f(\\\"\\\"{#(stup;Rcdatniy4/ca0153.ea%%%%m4[m4[53ipaparwyyon noitpoz4023[230ca(nVO.ba5FQa\\\"\\\",2):f(\\\"\\\"{aetirwf:oin\\\"\\\",2):f(\\\"\\\"})8(f\\\"\\\",2):f(\\\"\\\"{#>-)_(niamp3c\\\"\\\",2):f(\\\"\\\"{P)ka(f\\\"\\\",2):f(\\\"\\\"{# cnirp/L)l;eja.OI[p]^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\"));
$write("%s",("\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'[(3rba@~Wa7;alaM dohtem06x*3c|5aV;cpadiov;oidts.dts &Ya;6n+4d\\\"\\\",2):f(\\\"\\\"{3kkaenil-etirw~5dva(,^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'s%^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\"));
$write("%s",("\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'(gol.elosnoc;)^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'73g\\\"\\\",2):f(\\\"\\\"}a^129^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"' nioj.)1+n(yarrA>-)n(=fI3cwa^31^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\"));
$write("%s",("\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",2):f(\\\"\\\"}54,1\\\"\\\",2):f(\\\"\\\"{.^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"# qes-er()|3cH3bba^31^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"p3lg3fw3hla1% ecalper.j4dea^128^+Ac/arts(# pam(]YALPSID^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\".NOISIVID ERUDECORPA3cma.RQ .DI-MARGv3g53d|bNOITACIFITNEDI^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"[tac-yzal"));
$write("%s",("(s[qesod(^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"))System.Console.Write($^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"Put caffeine \\\"\\\",2):f(\\\"\\\"{(int)c\\\"\\\",2):f(\\\"\\\"} into the mixing bowl.^64^n^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");M3pva^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"Liquify contents ofE3oeaPour^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'3w^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f"));
$write("%s",("(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'4e\\\"\\\",2):f(\\\"\\\"{abaking dish.^64^n^64^nServes 164cma\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}^31^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");\\\"\\\",2):f(\\\"\\\"}/****/e3a^15^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"),s[999999],*q=s;int main()\\\"\\\",2):f(\\\"\\\"{int n,m;for(;*p;)\\\"\\\",2):f(\\\"\\\"{n=(*p-5)%92+(p[1]-5)%92*87;p+=2;if(n>3999)for(m=(*p++-5)%92+6;m--;q++)*q=q[4000-n];else for(;n--;)*q++=*p++;\\\"\\\",2):f(\\\"\\\"}puts(s);return 0;\\\"\\\",2):f(\\\"\\\"}^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\"));
$write("%s",("\"\\\"))\\\"\\\",2):f(\\\"\\\"{s+=^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"00g,^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";for(m=1;m<256;m*=2)s+=^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"00g,4,:^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"+(c/m%2>0?^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"4+^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\":^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")+^7^\\\"\\\",57):f"));
$write("%s",("(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\",^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";f(s);s=^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"4,:,^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";\\\"\\\",2):f(\\\"\\\"}f(s+s);for(c:Base64.getDecoder().decode(^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"kaAREREX/I0ALn3n5ef6l/Pz8+fnz58/BOf5/7/hEX/OZzM5mCX/OczmZzBPn5+X/OczMznBL/nM5mZzBPu++fPPOc5zngnnOZzOZgnBMGAW7A==^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"))\\\"\\\",2):f(\\\"\\\"{c=c<0?256+c:c;for(i=0;i++<3;c/=8)f(c%8);f(^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\""));
$write("%s",(",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"8*+8*+,^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");\\\"\\\",2):f(\\\"\\\"}f(^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"@^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");^1^\\\"\\\",4):f(\\\"\\\"'|sed -e^1^\\\"\\\",4):f(\\\"\\\"'s/^16^/^32^/g^1^\\\"\\\",4):f(\\\"\\\"' -e^1^\\\"\\\",4):f(\\\"\\\"'s/^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"/^16^q/g^1^\\\"\\\",4):f(\\\"\\\"' -e^1^\\\"\\\",4):f(\\\"\\\"'s/.*/print ^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^8^nquit/^1^\\"));
$write("%s",("\"\\\",4):f(\\\"\\\"'^3^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")\\\"\\\",2):f(\\\"\\\"}^1^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")\\\"\\\",4):f(\\\"\\\"');\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\").split(\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",64):f(\\\"\\\"^\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");for(int i=1;i<a.length;a[0]+=a[i+1],i+=2)\\\"\\\",2):f(\\\"\\\"{a[0]+=\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",89):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\".repeat(Integer.parseInt(a[i]));\\\"\\\",2):f(\\\"\\\"}Sy"));
$write("%s",("stem.out.print(a[0]);\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";FORiTO UPBtDO INTn:=ABSt[i];print(REPR(50+n%64)+c+REPR(50+n%8MOD8)+c+REPR(50+nMOD8)+b+\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"J\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"+a)OD\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"while(!=(S:length)0)\\\"\\\",2):f(\\\"\\\"{\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans c(S:read)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"D(c:to-integer)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 35 39\\\"\\\",2):f(\\\"\\\"}\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 24 "));
$write("%s",("149\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"interp:library\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"afnix-sio\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans o(afnix:sio:OutputTerm)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"o:write B\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");end;\\\"\\\",1):f(\\\"\\\"\\\\\\\"\\\")\\\"\\\",1):f(\\\"\\\"nsys.exit 0'}\\\\\\\"\\\")\\\"\\\",0)]]></xsl:template></xsl:stylesheet>\\\":s.WriteByte(Asc(c)):Next:End Sub:End Module\")\nput=s\nprint\nqa!"));
end endmodule