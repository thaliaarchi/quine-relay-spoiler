module QR;initial begin $write("%s",("Module QR:Sub Main():Dim s,n,i,c As Object:n=Chr(10):For Each c in\"<?xml version='1.0'?><?xml-stylesheet type='text/xsl'href='QR.xslt'?><xsl:stylesheet version='1.0' xmlns:xsl='http://www.w3.org/1999/XSL/Transform'><xsl:output method='text'/><xsl:template match='/'><![CDATA[write,format=\"\"%s%s%s\"\",\"& VbLf &\"(\"\"\\\\write{-}{txt}{(\\\"\"with Ada.Text_Io;procedure qr is begin Ada.Text_Io.Put_Line(\\\\\\\\\\\"\"print\\\\\\\\\\\"\"\\\\\\\\\\\"\"STRINGz:=REPR226+REPR153,a:=z+REPR166,b:=a+\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"2\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"+z+REPR160,c:=b+\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"8\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"+z+REPR165,t:=\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"write('implement main0()=print(\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"BEGIN\\\\{s=(\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"#include<stdio.h>\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\nchar*p=(\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"Ra#include<iostream>!nint main()\\\\{std::cout<<(!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"class Program\\\\{public static void M83abbSystem.Console.Write(!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"Quine Relay Coffee.!!!!n!!!!nIngredients.!!!!n!!!\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\");for(int i=9;i++<126;)[3pva$!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\{i\\\\} g caffeine \\\\{i\\\\}I3b54rja!!!!nMethodv4f\\\\{aeach(char c in(!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\")))s!!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\" [2b.a!!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"rts(nltnirp(])]!!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\".NUR POTS!!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"!!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\".h3bca!! h3dA3bha[))!!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"e3aea!!!!!!!!h3d[2cga\\\\};)06xm3f$3lpa)1(f\\\\{#qp]\\\\}\\\\};)0,#3rv3rR3sv3mba323284-fa(f;)1q5.ba.>4[ga#(f;)3P6[=43ba7=4.<4[<4[<4[v3g2=d=4[=4,kaD ; EYB RCH4[H44da,43?4[?43daDNE%6[%6[?4;ba6p=Wj4d1E/*D[*Dbca Ae<[>8[?4[v3neaPOTS&6[&6[?4[K9oJ9[\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'6[?4[v3loaRQ margorp dne06[06[?4[v3kbaSR9[%6[?4[7P[\\\\}6[?4Lba5/G/=4[~6[~6[v3kba&f=[$6[$6[-@neaPOOLwN[,6[?4[v3nea\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'&,)&6[&6[?4[wNmga. TNUON9[+6[?4[73mearahcE@[(6[?4[P9ngaB OD 0zN[,6[?4[7Gn33)>4[#6[7GBca)At=[&6[&6[ZJoUJ[\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'6[?4[v3mqaEUNITNOC      0126[26[?4[pDmT9[%6[?4[iDnD@[&6[?4[C@rba.(6[(6[?4[?4lja1=I 01 OD,6[,6[?4[?@meaA PU)6[)6[?4[v39<4[\\\\}6[(NBxa;TIUQ;)s(maertSesolC;))T4[96[?4:ca13@4.banl41ba2l4/07[07[?4;ca36#6[#6[#6[?"));
$write("%s",("4kba20>/ca\\\\};&6[&6[RA<ca52A4.damif(6[(6[AA=ca15@H[#6[#6[H9?ba+E9[%6[%6[v3m%a315133A71/129@31916G21661421553/c5[C6[C6[93meat+s+C4[(6[(6[S@[#6[xD[93~oaamirpmi oicDAx\\\\{41ba6M>1baCo42ca779M/l41ba0j4[ga#(f;)9-9/pani;RQ omtirogla99[z;[>>[hBn~anirP.F;\\\\})1+69%%))n(tni-i+512(Q3)C6[C6[C6Cbaw?4[$6[$6[i:nhaaepeR.SwI[-6[-6[v3mbaW?4[$6[$6[v3lea=+s\\\\{tW[(6[(6[v3m$6[$6[gP[$6[$6[?4Mda320XP/da\\\\}\\\\};(6[(6[?4;ca40I9/%T[j47da345@8/dadneA8[A8[QB=ca62RB/B8[j48ca38B8/naPUEVIGESAELPnz41da289z4/76[j47da411P8/ja1,TUODAER:6aD:[)<[lB;ca86L8[L8[tKiba4SX0\\\\}aetirw;\\\\};u=:c;))652%%)u-c((||z7[Z8[5K;ca73Z8[Z8[jAhca27Z8/da#-<[6[@8[?4:ca88wQ0@8[j47ea7003m4.da||i(>[B8[$Z=ca0867[A8[@Fgca92A8/ia#BUS1,ODd7[D8[D8;ba1\\\\{Y[D8[*Liba5D8/mJbia)3/4%%i(|41qW[86[.Yjca2886/x5[x58ba4k4.ba)M<[2>[?4;ca6"));
$write("%s",("7<8[<8[yLhxD0)[[B8[?4@da974B8[B8[UBhca16([6Na2=:/t;2%%t+2*u=:u\\\\{od7 ot0 yreve;i-=:u;1=:+i\\\\{od))1(evom(dro=:t elihw?s;)s*9P[89[?4<da41189[89[mMhca899P/ca-<8P[C8[?4>da528[L[C8[j4hda7219P6e7[E8[E8;ca35E8[E8[j4hca65E8/banVA2sV[+6[j4ida238+6/ladohtem dne.662da189y4/66[1W8ca11O8/ganruter162da30716[16[x5hca9316/CaV);gnirtS/gnal/avajL(nltnirp/maertStnirP/oi/avaj lautrivekovnin72da963n7[n7[BEhca275@X\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'G[\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'G[sWnca80=8[=8[+OjpU[x5[j4hca82x5/eb\\\\}\\\\}\\\\}\\\\};0=q;)]q[c=z(tnirp.tuo.metsyS;)0(tArahc.y+z=]++n[c;y:]q[c?n<q=y\\\\{)0>2%%++i(fi;48%%)31-)i:3c&as(+87*q=q\\\\{);62061<i;(rof;n)rahc(+G:[,<[?4:da104c9[n:[+<[x5[x5[x5[x5[x5[x5[x5[4VGca86vK[HA[HA[HAjca31<8[<8[U:[x5[x5[x5[x5[x5[HW9ca77\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'T/oa=]n[c);621<n++;Naqa0=q,0=n,0=i tni;u>"));
$write("%s",("[U?[?4:da0006[Xf9[#;[x5[x5[x5[x5[x5[j4;da809l</$b6aeeicpbocKhLf@v6gX96gt|\\\\}bJaMa\\\\}bJaPa6gPXJaJaUa-bJaJaTaJa8bhw;a8bHwKa8bHwZ=6g+EOaSa;OFHKa8b;ON/8bGvHw8b@v,EJaLaJa8bGv@vj4coa8bNa>|@v:b+bX9(4aia\\\\}bJaHaJa93c>bHaJaJaQaP0;a8b>O:aUa:ahwocXbddxepgXcVcScQc/aDg|bjwIcncDcaj@c|bKa<c=a0co52a;c9c7c6c4c|0hN=aJa|bxekcpbzc-bCdlepbocHazcHapb6a6aIc7e=a-axjed3bHd6a6ao3ada|b9i3fra:e7apbk<FeDeBe@e9m3dEa/hjdif/b/gdg3fM+zb7ak<-h+hMaxjed-eY\\\\{Ja>a2a,g*g|hMaxj|bCfXbybvd6a13i8bHdGZvdie=aSexvOa-axvOaX2gbzuSe@hqe7b5aIgjcYcWc6aSd1bji7*-bChMbUfUfIb/bHdlfjfug-b1bQzHd6aSd?bpdX\\\\{n99ati6aVj2a5arifeefdcNh4ajcJg|b7,jc?a>f?h|6ak3aeasi<bx6albkf8hNdoi1B:ZBb@b6.;a,bpid*fbpbUrEU>b37PfLYyg-avfP\\\\{>f3hCd1h:gEaAe4gyhwhSf9a7btd-a5buZ-bwh3a=a9a7bp@s3g53ecawh53kG3a33iha,b9a7bn[3hyaFa>,Kh9aq-xb-ap"));
$write("%s",("JXklhvg7h\\\\}3ak3asaLi=ekfwh3asbxhEa3a[5ak5auaLgxhCaRf6a@h>gOgLh:gk3ckaVhuh<b3c-ao7c=3geaBeRfB6ao3aja=h;h6a<bxK?[v3a#afig*oKb2a=lSgQh8fwbXcjc@aCcVc6.>b&aub5c5aye=anbSgybph5a\\\\{e6a7bJgHawbXx<bsa-b9a9b9adhSg-a6a>ao3aea@a@aq3a)a@a0c|b9a0b9a@a>a7a6a@a>aIa|b>d9bJa0b-3a%a-b9adh9aCaAaJa9bSgnbJa6a|b5a,bHaJ4aga-h2y-aa=a\\\\}aFt/fFt/f6a8b5agq*e-a=lkLbb-aw3aba7w3jka=ljdEfs1Hdx4awa8b9a7b5aMaJayb>aoqGa1ci?awaHajgJa,b5f1cJa-b-a\\\\}c\\\\{co5a%a<aSdW9Md:aKhJaub.e3fP\\\\{7*-bJa3bjce9cgaJh3a3b2<e>8aDfUhSh;aYcWc=lG*,eJi:i2jnkziijXj*czjskbkChtF4qVzuboYT-;mF2+-Gai2SaXk9<@?O0g1:@WC.bTaxfe-CaW*BrZaWnL3lb.b6@WnYamu2@-bV<f8Uu.l8Ldbt\\\\{dlBaZahbdljbIt8Phb@aTaO2Aa6oYaos@oDaY\\\\{mNFhibCavMI+EafO>\\\\{>aYa0wMp>/6<W0U0s2vbO-cLcbvOyo-\\\\{K7k|3lvb*/>te\\\\{>s\\\\{byF8Qi.+lBvaofxmb:0YaDr=aBa2S=aV.WafbZaV"));
$write("%s",("w+b>aR|xM-b=a?VFxom\\\\{PnMkE3bU.\\\\}<ab;*,Mbom+rwSu*lk\\\\}Fxfbl/St8bj8HRP2.bbA/y2zbEiV/PBjdbHsEn*bCltRUhBejb,bTazbp;\\\\{:pzFse5r?>oy=4rl6Wtg1oYiojbet;k=vxOnl5b:>x@AZjbeGYoFae1TaAag+fu?/ibWa3zb4Jp/qx\\\\{I0SqV/XtRlhbndmuOagmgbg/.QSaBafu.b4sTl>S[#U[?4:ca36@4.ia(ntnirpns41ba2AO/ba)R5[77[77[v3kXdI0EwI00pXa:AFx1m\\\\}EegzmcmOaP2G*yb=ahbvbgbwyabb+nn.b*blOkbWajPBa:U?tCaub2gCaLp6P+mpN57EaP2G1CagbvFgJD=@atbos<aubctEebbv;UvJ8VtFufbFawA\\\\{bPQOIEaxp4k5bDa-bc32b|Sc|TaR?|Se-8bZa=A\\\\}vMsJr9vTa6R.kBD\\\\{dGkCkDaPa??I94Dh=WMcbfbC76R+-G<mbjbDa2Rww7*\\\\{bSa\\\\}.F8Aox?6,u?abAq>aq?z*j:y\\\\}l?j?nfh?f?kwjbDaO,2zQ,\\\\}.SXjbDaTa?\\\\}Taww\\\\}.3bWaw\\\\{\\\\}\\\\}4zApQxC\\\\}.n/rGySr,k-lG*YajbMpDaMc8Lc3ckcQkUa*P2>Gywvk<by9>NrNRgvwHYp6mQ,\\\\}>Na2kOGD*yzQDilUkGy=k@nR2E?NwNp@v+n.kG>.kplvb4k|x|S|g+sA;.\\\\{A;+?H"));
$write("%s",("wxfNJ\\\\}.9bRa+bGyK9GaD=SaUu/k7lnf==A;:=A5xA*v3IBmDa9bBwYaosuudb/=7x8Ljb.b?aebWnkbDajb.bTqk3aHb6d8LibAab60:*y0:*mdbJd0nG,8P+,YadbEa,bcb7?EnI6hAjb.bWqhb2bz<OM?@QkdCe\\\\}\\\\{wV77u4wCM1|.Q7b\\\\}khb2u:81leli9O8H<F<DTC<1lcn8LUFbs,k@9Dasve\\\\}:s>a.bhb2bq<hbpK>n?ajbNaq3c\\\\{aNae\\\\}c\\\\{Gp4qhwhbNa0.0bmbN-I>)3e:dEkN-Bx=mhbTlcw1lPa*n>a*pAaBaDa:sHtub?aN>U;E8vo>AEa+mjbvoIkcb@a?->rY|kbab;k9bw02bowP*@amb2bZaFaQlOl8;XaNp5;3;TLwbprSa2bpru3+Evb?rD9SavbQkA>:85L5eMSK8mD60LU9zD5mbX5:AAa\\\\}tvb=a@aL6jUeb6b1b\\\\{>J3ib-k|wN-wy-Fl/B\\\\{-bBTXahb4A+wBeYl2b10fHTa60KrO8F<jov0T57b.pEk=a4yfzk\\\\{1l>nYaYa8Z8bDa0b9ze\\\\{C7qw1HMS9-+bYaibXaJI<-*0/C.|kWPrgb\\\\{wfb%3[<lRam:3lly/yNz,8Wq:v2>@a\\\\}AhpZymb7*Mk1+DkHfhN\\\\{ZuUN;tb\\\\}.>,Bak\\\\}2\\\\{dbBgurBg|lI<hN1c+bb\\\\}G*Jrpx:xjbZnO86pZ=qDL8YaQtG\\\\{xfYBV.zb0<=tct"));
$write("%s",("dw,8I|wdN|8c\\\\}bxbmbLdbbF|<e*;cp+F5FvddbQ\\\\{\\\\}S;F6bI1lb--wzl,A?VX|,Mru?T:jJglzb5bStjndg6qH@Xaz2\\\\}.GxCamn2Dcs=*J,YaYar*otOHXkt9wbdM2bDGm;Auq/S|prBT2tR19=sqSaH;4Tbbg32bCaNaXt?aRtg+Y3Aae:.u5bbbebab1Bh4o2z8wx\\\\{kL++eg*EDYpF=AaZa8uorRoAudwbwvT>a*?a=C7QVTST71+dt8beE:A|9Twx+A\\\\}\\\\}b,bvuIN9pus4bNaPBZwtnXaUad<*+2\\\\{Vad<HvCvtq*bip6b6\\\\}|c7vHx@?I6?-uo*bIE-Z=v;vvz*bD?lxwp|9af+EgMil3l/yA5yREylq=AV0EpyPf1syBDDaOUQ*.p7b5r\\\\}b4bdb7Nk*|Ig/Bac6nw2s>|DRLylyA,,+Uajb0|IqDRWn/-5umWyuUagb,yPwNw<NowRm+zL@ow|J,zgb0uh2R|Fa+IjwPaA1,EubZoQa6bjJlq;I7kibgy@XWmUy\\\\{bG*0<R4VtPnrVNnYmub7zsukfKL*@PkfJty0z85FxV\\\\}b4av=hOatRAL-sI07+.bX076Fas6.4?-4rybBvp5D|1XRL:A15n66z60,s@nZaNrluAvcN4sIkWa8:?3Va>aG\\\\}yRSambNr3bK7fNAy\\\\}QXt1v48\\\\{|Qaab@avbPSe@\\\\}S;Fb2v34lX<t\\\\{ybhIp/FsCTtv7*5k4=>Ljw5kubgjo"));
$write("%s",("vEnT0EDgot\\\\}xpSXEaPy,eXPWyR-kAubYMc;-wW|\\\\}Y9bXa,q-yz+@XGDwbA8Qa;*jAftwbLIx5Oat+5\\\\{OaEa.-pqBaQ|mp.==IU2WF;xWa;rQa+jOkD2XoEalbfby17K9Xlbg54GRaphNQ4bOa1v\\\\}bhb*xybbo**-3agaibsY;x\\\\{3a+a22D3/bO,OawbGld*.bGaxChbLu|w,b?GboRpEau3ahgboSn/M?=vbJ2\\\\}b|3Oa.HO,|bOakbRuAaj9xkQ4ClB@ukvyib\\\\{bj/l<ftXaeQ:8BAzb|ZpZy+NncmphOaybkbWa>a2ylq6nKPH@hw:Dzde-e\\\\}8vFa@b\\\\{bF|rK8bUKPl2yjq+pO?bbu6Xaybswbuvdn6xZ|0\\\\}dVa?aQ5*b=a7s:zJ*F\\\\}-bH0mU,*e1wq|y:Dur.boZ?v4bAaO8,bhZhbNf@nDacb|.C\\\\}g5ag1,4vYa:xI?PY+wL6llK9BD|OfAao6b1r3COHU@*u99NaB>O||b2,V3+bibZa+pflvwZng.abI1K6QRLPY:Z=F8KPl6urA-jxrxAAFaNx-\\\\{9bDmY?/n?aubFaz4,d49Uu\\\\{bIy>0D,Jmcb6bdbJ:Xa1bCrAvpH40Sq>7/:I0\\\\}KVz0IOLFrS/8UOWG0wb\\\\}.,C2bx+b8-b2bSu-8:mEDG*6wR4.0R,xbOrJsYa@5eba<g7P*9U-bvO.bHt75lCtbD3NOS+2bpJ\\\\}vdm2sSpJ1-bu51\\\\}.\\\\{plu"));
$write("%s",("fa8\\\\}brrk?d2Kn6q,/82PCS1ba0BS.c1sfr|b8R*pVqe@eGUpTTA>.pNaxJ,:Zy.rkbAOX2bpPaG1E9c6NfsS7KuOW46bnqZy?Ko/nqLu6.dodPUh+w4A=7zt=7I/6KF<lMVaYao@I\\\\{+,4/v;*J+W@Kd4hI-b-9+bbuNa|Od4R,Jy?qd4?a7\\\\{;S71G|DangYps46bNaK:/\\\\{??L//bibG*,b7\\\\{6EUH2;D0b6z4BaZAP*Qa-\\\\{;tFkYa=7cND;zborWsb6|gI?;DEnM6YFDa=a23\\\\{bjbz\\\\{?7Rm2gtsJuL3J.DK:uuq;4b/;nFyjb*p<Ihfh204.4xJBaLqEUT5ayxf<2PsuqWa=7t2-bO8ubuOLey+6xkrwb0Khq4v>*Z/\\\\}bbteb@\\\\{Q\\\\{,7vKqvFa.uJte\\\\{@50p7sV0MqG11b1@Ra\\\\{s*@EmAaUa6./bm1Fa6mhllC;vGf7rWs8;5b?s5nuy\\\\{rJ.,p\\\\}.R20y1CWa9\\\\{4nDqlxjb6lG*q4>an:XkMd7ln:loOazqBf;z4f@l/M9wGN;zGaoKQLxsrqpq,bkAEaKdiq-wN<jsCaL5XmEeGNuxzJ>ejoWaYa*/P0xbVus|z\\\\}\\\\}A|cN<\"\"),\"& VbLf &\"(\"\"yb?3Wm1q<aiG;Lb|/|gb@a>3kATtg*Q|.bO|rIvAcwC24b9@>K6bzkcsBL=pM7Ga>8CtZwkAYpX\\\\{R\\\\}6Oo+3bJ2IwcoS\\\\}7mphqDwktby\\\\{,bPk"));
$write("%s",("ubNFFnYaDpuB\\\\{bPv3QRtC2g-YazuCkCa\\\\{kkn?a4I=o1b7L.bYa\\\\{@Yo=o=EX</bYaFahQ60G*TshNVPBaEa2y\\\\{O*v*b.nN/mxlCjbZA@apAA1?sSlgoRBQ0T:Som0/bFke@8*3lZu3b|86b?ayb9bW.Ly*-xfMmyFSabbxb441b7wmyI?-b*bZa-nO7Qa=PibTr4shyVz:7VaPaALlb?30zu./?D-mR:N\\\\{xu5Vaq\\\\}Pp:uu.b3\\\\}E|bA\\\\}Eslir7,b..q\\\\}6DFL1k?kRHSaQxPQI1G|Y1SGu5lbo+\\\\{/+k0o4OXtVt.-qPfbmb>?tbzbmpUamtVaHlDO7\\\\{H-E|F\\\\}:?g>b6vb.QUhCa.-Jrptvzcb7\\\\{G*RHGAmu:kxfbO/@z2qo*bc\\\\{ZNCpXt6OMvsqo+7bbC6|=.*l?-G\\\\{9t0OvAl5nC7+09vrKsks|bJ8BFBa-/hxgn*JybBatbY,Zafbp/604zQ0m1TeB1q>@aao3b<albif+?Nw\\\\{bzbe\\\\{UhL|YaX0Z;J?Oztpb+2bcJ3b,lEfQybbZa=9mbauSa-5o2-b:pUy+b/@ibkfd*,EVs7?*F>aybDm9lk*lt>a0b2zvr5b7rgATatsO0myIt\\\\}?0;w8i\\\\{+mW/GaU/nEWa=\\\\}Emxb|bCa/bprg*LJg6DLVaWau;M\\\\}ebG*@\\\\}UaAa@\\\\}NaG,zbbOc.Wa7bryG,B@ONWaMNa8JNHNU8Va=iT0abH0b5/bM5/b/"));
$write("%s",("b4r@oh2/mfOeC?ao+lbMq?a7AtvjwDac./bGN*bVqyBEaTan7pp8t,:Ct/bvbAaOavyAa+b61dbjbVa+bEmw1-faox>Anlyw|?q;n\\\\}bmbW*vFkb3s0tinOJIdKd@?jhsrG|5\\\\}|bTag\\\\}EeO/-@+lUE6\\\\}dM?nQuD4vq9bNaYazd1C@ab+vDDAUhGaX,?\\\\}ubiFhbUaybG?Za<a,b.2?q\\\\}E>m88\\\\{-XmBop2>a6<OxUur5lENrd2vbFtHKLbW:/xB3fv*bCoe\\\\},bbA;zO;dv*-K8M;3vVmB+0bE-yL0k<+>s1?xfYt,8oy,qz62b0wOaD.vFd|<C2*Ya|JwbiDjvEnblUaYa+b\\\\{bG+9b2bBaQaJdWJm|nw,bVajb0b1Hcbg\\\\}yHJs5b+Dx+H5=a/b\\\\}bxfuG2bFaV4J*+bu5Poab>nAaYa..J8gbZaOaFaEa.\\\\{t29Bs@ctHCCtxfD2<e7K@\\\\{u3Fl0*ag0b9=fb\\\\{rdhlLHAGaNm.bp|*bP2Jl>rxbjl1b-9?KJs<KcbP,jq5bPsoxh|zbLm|n?q7b8K6Ko;=lS9MG;Ipv-b44+D?qLDOaPani=v4I7rj6*ycbwb>7\\\\}5=v6baxT-\\\\{webCa>e.qP6CaXav;Ao;r@vafkb/b-J,7CamKxfOacb.brJ<arJ?aSa3JctO9D|hbtb|bu5Qpu5fbCahzY9=J=Izn@J1bSa|c.p5oMs53N;mb4bibQz7Jhzi9mbzn1s5\\\\{uJWC1J"));
$write("%s",("tt,7JvmbQ-\\\\}JcbI<XavJ-J:2tJAf,qzbV\\\\}ebmm\\\\}br-zb1k3bsycb\\\\{62;5b.b1k@alFTaTrubk*?@Ga4uhbIshbjhSa=acsDapt\\\\{b/CfvVt+IfbLl1bzur-G*+,xbabts@I+,xxRa5bgpOa1b2yjylbAv?aBa@5JthlT0iDEaib\\\\}.D|Zav@W4x1WoPaly7sD|,1Zy7b\\\\};*-p>rt1b-\\\\{abxrgIjbZeC2EBindHD;<aVtN>zd<awbYpo/Oafbg/XnA4xfSGQGTa2y.-ib=vXaGw<|z\\\\{/|.\\\\}x\\\\{9bab75+76\\\\}h9v7Jt6.UaS4Aa-2\\\\{oNr0/h=\\\\{b=alb7gabdbEEWaBajo*F85b|@?P*Dm?alb2bWajlklRaBa5<<a>>A?\\\\{1KATmNajb?az><aNrfbjq,E2gllCr*GQpow:2PaWakbnuEaVaG*tbmq92-lT1W45j|AouSaOtk<3mX0\\\\}bybabQ.Z-Za>bblZ01bwmlbBDfbc6Q6f.Gxg**2j@/0;rU.m|mq8l+p:?jwgbe,\\\\{b*0g5Sa9-@uRl*b>*Gal>NwUkWaCaC2tbl|wyfw5,B\\\\{tbabhbRwR40|>vL\\\\}J?tbJFurtb6bgnD*M+D*e@C/9*tbFa3z\\\\{ktleb6-QazbApvd>vx?:/bCT;tbXoAowbqmDag-*bdb?ai:4=P\\\\{kb5lb@ebP,bblvOtZ@or/b28k|XaowM6/bnf0+ubBa-bCaBfBEkENaFEXa>"));
$write("%s",("<E1ubG*jbW\\\\{Eu@7gb7dpo,EcbTas2JqDatbo-mt:E:575/bEqCa>jeb4bgbq7nplpYqubqoF=ibDaVarq/3\\\\}bPa-f\\\\{byb/CYocb5bfvZuzbv>w\\\\{ab4dL85.5bbCgbFatb;sd=TaLvYaZ0Nl5b.w\\\\}qC\\\\}J.xbyoqqu?ybhbfb8bzrebG4/bb6;*7nXtpAAl8b82ws\\\\{bu5?=/|xo1b\\\\}8zbvbMo;rTp8bM\\\\}>aYBur\\\\}5tx;rjsDlebxf6g,mzbD0/y20QafDGaduu5;mfv8b3tEzzbZa40z4ulcbu5/yN2Auv;*;p;O2ouQujplbZu=9G*x+jlms7wDCXvKpdq\\\\}:7?q69bxbfvc//pvn|bnCftAoYbTafbgbItRaIoXawp+?mn,7IzjbU3eb=48y,pMlUni6abK8Svxf2bpAQt@\\\\{4fA5G4ibV7J:0b5r.bB\\\\{Cr?a;qRa\\\\{b*b:2VzVa*18:@aabc/lyqAb3x*\\\\}tr5YaI+fktpXa=4Fas;9@KAQwNaH5-4Oa\\\\{1:sx+l</linN0=\\\\{;=f8Y<bp>a-bDaSrxfwm1b8bNf>?KfJr?-0<Ct71+begYa9ohbFagjJ8Zu99S@6bEaAjx@@50byyvs9bjbU2exG*Ga14w9@m,bQ4>a<+Aawy-wPmQtsvVztb<aioN0Oalb|dgm6bOaDqybhmUrzqOa,vomyb9zH0DappO;Ua*AKru33lXr7b+r+=Kh|bZa>a2z;xGaRcab-bSn"));
$write("%s",("Qnpx=a-bXa85jbRaXuibZyrx*b0bVab\\\\}4bmbXag>/b\\\\}.cgTwAhxb+5ez7b>-q<-tL@<@\\\\}bWsOabbtbr\\\\}PrL3o=89Va>v<vabOtzr89FrjbxbRa1vZaBpnu+t6yQadbkbu4?as@A;3bGzG/5bPvX9RaAp2bUab?PaFnubxbT.Hxu\\\\}HvCrGat:zdZ9l\\\\{lbwkhzlbGq1b1b91ao+tQ4mx21O;KijbQaz<G15oe>>aOao05oV9cb,b7oybPa!!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"!![2fha\\\\})1(f\\\\{#v3rga(f;)0,73-c1wbTaRamnJ88b7bOxfbXaql\\\\{m7npt0bvbhy@\\\\}xbtb@akbyb1bKi-b?7wm/bGpvo1b*pB>Wa=aSaC\\\\}Mz90zbhbur>=7mzbLke>0\\\\{?a3b2z5qg3+7\\\\{12t;\\\\}Gok\\\\{-0t+UpjbubHdB==ah0=aRpkb6-wm<>:xDaNafbWtYajwg*Kfn1*z89c6AgwrNr8c,bG=HqlbT2abWqwvt;Sr\\\\}r|b,b\\\\{tRacs\\\\}b?aQwp2tx\\\\}bNatbOo?8Fajv+1Ua6b-bXo,b;ryhU50oTaerG*bbjbRwy4dq6=TaD*>0db"));
$write("%s",("+19bVaSyXvcsRa0b@p\\\\{b6-Mlw9Fa2b3t.\\\\{w90b5b@a@5z289+x4b9b-=Naj-;r2b4.ru=aNpJ.Ba>kZwZa?vo2b\\\\{o2v.61,*b6Wa4bg*\\\\}b1su/NaJ*Xam|z/p/xbxbFa1g2tdbebt|>7k|g7x7psN<ni\\\\}b=a-wwkybK+wb|qib0bHnlq:<oucnAaP/v<Z;ubhs@blhZt3:kb*bmtf|W*=uxfA+>jNar<1-4bCanmitdb?-+binablpN\\\\}E71s\\\\}b/bTaXaavEa|bgbJ:Jp|8-bQr4bP2Zu-b6bG*+1ubm5WbOa:7n7bmwbRazb4bI0ptsqGvgnJkU+:;zb3s/;jb-;Ks-26\\\\}SaL\\\\}/n8sUaSl9tm0RaqtQaR/Rary8lXaLl8bvb+b,b/,zb946bprWalb9bzbfb,wubEa\\\\{bVaeg1\\\\}q6+m\\\\}m\\\\{m9-=azb0b;ndbj/P6PlV+Hu:8cbY\\\\{Lud\\\\{ib2b9u=u=9zbWaSt460|p5=94.0b|-q6|+jobbNc3lNvLvZmwbP\\\\{?yMsi:Ta*eAm+bwbcbC\\\\}bbAu@3>agb8bGrttJqvb5\\\\}xfxp9b3bebA5Zn6b/bQaTajb>aCeO15b\\\\{bRpO87z|yGa9\\\\}+b|bAn4w+oFtazPmbbQa5v7o?bkb1oPaQa\\\\}3ffG4|bYus1ArPaxfRwgbw9@o\\\\}kBalbXjH0tdlb@ogzezjb*l,pjb4bv+Ra|c4bS\\\\{Sa=qI8wbg2FlAaGpu"));
$write("%s",("6NaVt4bybr/g/71NaCa.bai<-q+lbdqhb,8T1tb136vf/5bkbjwE1jbCe.b25=atbwbAa=aR.\\\\}4OaIl5yN-Kf0bk+xf8k.bcb-|*bmbub<|=*g,mbo|m|N1zlAxH5tbxftmgs8bmb9ujbh|T0OaYmKoQkXbt-Wo3dL/HnNn,qU.ubw\\\\{w\\\\{2dSahb+5\\\\{x+b@ayb?ay\\\\{oqcbOsG*XnDv1bjv4b0s<a0tZaubvu8uAe\\\\{bin?sXawwAnOaYaQa2bM6>uWa@ad.6\\\\{s*/b.3,bBa0z;.U+\\\\}59tUabbTawy*bh23dlv0b:sEa<a5bWvbbgb3bs\\\\}PaVnTnNcvb<vTl*b41p2byAf=u9*t3mb7m:d=piuk\\\\}FaL*3tbbXaJ,DaybJ,X\\\\{vbD6BeAoPkS\\\\{@qDadb<+hpdgt/;mV..bVq4y0b4r6gBa7+?sv6t6<ointl/bP2lus1lbwbfbQ.xz3b.beb*bVa>mTaDaf5vbbb8bc\\\\}.b=u>ngbU5>a7g?afbAu9*go0b\\\\{5Stfb*bEaq4G*v\\\\}Q,Dahlxbp+.\\\\{\\\\}r0b|bbt-4hbWq.uUaxf2q1kxbou+1tbj/xbhbUm2b7z@m<aUaI|Fo9-ibVv5b4b+bbbZnW*qm.b/n/bUaRaAvyb\\\\}q@aEahm7bZwT2Zwf5J4\\\\}bOaBa+1<aQ*rp40Ozq42bdbgbQrzb>aPa|pomwmbuibkucb+rRpjb=a/yibg+Jp+bom5\\\\}Cl6b3bMqrs"));
$write("%s",("YaGhSrL|Vmdbzrgm|b<a?aFa7baf0kwwYcg\\\\{8yvbCayblbtbCa2sRa4lOaTa6bql,.b0119rh|kbmt3,<qebtlTaF|,lib.-1,-\\\\{gbc34bfbkb9br,P/K*Ea*sG*<aCaOa7bUr?aWa\\\\}b6mmb8bib3dGx+p;dnuUavwFxS\\\\{\\\\{,Z.yb6bpowb7zD+|bIn\\\\{z*btb\\\\{00b/b4-r*Fa5bvbUhjtxx5\\\\}vb-\\\\}ZpprZ..n7\\\\{x*\\\\{b,l*\\\\{Zx7bbbe,vbW*Ua,bc,|bVablNa,pZaibTa|p*b>,VaJy8bGaLojoebibwbBawb;.x+FvOaXmAa9bwbBnbg.wZwhb?a1b\\\\}bEw6bZaAq4bzb1bGq\\\\{rlbW*4bZ0\\\\{bgo?aXangAoubYaS\\\\{2slxXcV/jbmb0b>/Q,UaRn0bbbo-xbcbtb@zZkUa1bZawyHn8bj|>/ct9bPaCaTk+b>j8bFagsUa=aebQa*\\\\{FangTahbG*Xa@aVa,,.bfbtbcbE-ybnm<sub5b,b7sy1xf+\\\\{ib5bxf/b@aW\\\\{/bBe?b5.80Na-by+ilK0cbEz,bFlNa4nppq|N00bOrOa8b2bkbmbu.40+bVaUaNa.uA0@0W.Fa0b*blyp/\\\\{b4lUnGaxfO+\\\\{b:xWa\\\\{||bNa/bFakb<hOap/OaNaxfdbc|tb?qx/ub@uGao\\\\}XrM/=\\\\}EaYay/9|DntbTaZ,lbQaFaMkip,bs\\\\}Rwn.\\\\{tJ.zuAzWaG"));
$write("%s",("a<*|q*lmbxfUaBj|.\\\\{bYaab?aTa5blbq/+pNaZaCawbqn;nAaowfu7pg\\\\}OaymW|>s1b4b\\\\}vWa1bNplbxbkbPombFaG|xb.bdbwb9t|ktbeb.bwyG*Hn5bPalt-b+b2bVa=ktz\\\\{b,+kbBa/|mbu\\\\{Pa*\\\\{yb+bpqtboqzbTaibOa\\\\},Ju=abbxfZnt-6bQa7w0bDn-bwmZwG,NkLkWatbHk6kWaSakz=aOaJ\\\\{;qjxPa3bAa\\\\}nmbP\\\\{DaEffbOat-lbipFa,bInX*\\\\{bmpq.3b@a7b\\\\{-Ua:uSasukbT->jy*4kCa/z2bibUa>aWaPaiwmbB-lhRasuVt5b2bYaRacbBaab6l*b7lPk@aWaww,zdb@aqo>amt4-\\\\{b-btb7bl\\\\}hm=adbrs3bKs8bMr\\\\}b9bAblbcbFnDp,bDaAm4btb|,Aa\\\\{vDacm7\\\\{gbbb7bwbZkmbqmxyubfb=a*b0tjb>pDahbLnG*=a\\\\{bxfQabt2yEaPq?aPaEaXaOaW+U+Yhdm+b\\\\}l4qWaoz2b0bnv*l8b*bFaCaVe?lFubnmu4b0bUp3bltUmYwwbwb*bfb.+hbCaPaabbb.bt\\\\}@a6g\\\\}k*bhzTuPyb|Z\\\\{yyct|b\\\\{mNaRavb1q6p|p\\\\{bZa*wcb7lNo@oN+oycbbbFazbUa3bN+=*lb3bxbgb.bwrdbsrZabbYa<adbabibTlGafmibjbMu0|*v2bRazy;mnm3bb\\\\}zb7b1p/p"));
$write("%s",("s\\\\}Ba7pDvev\\\\}budGamllb+*vbHlAawl0x3bkbTaZ\\\\{ibwl<a;rgb/bRaur<egmNaPa4s+bmbbbkb*l6k\\\\{bz|W\\\\{ib,bLdDaGaCwkbFa;k4a2|S\\\\}3tBaNrBaau,b-lxbxfvbZaEakb,b4bOncbFa8kvbmy6b9lYp3bhbcbRaTecoL\\\\}ValbNa>mUarv8tvwWaTa@aouHwWa;\\\\}Aa:vXv+jkbyu7z8bftSaEa/bktOpCoQa0zMelynnD|ktNxWaEaSaqoE|C\\\\}ty.bRavwVaTaIyVaSa@aNx|bFxSaxf3bNolyNa1b2nWa<w\\\\}bwsylcbDaSaKp>p7g4bdtnm|bRa=h.bWaZaabOaAaxfubTh0|kbzb?lw\\\\{lp5b:uDaszTaab9bCaibqq3bnugoCakb|bQa|cwbzbEzxf-bkb0bgoUaPa7bVatl*bBa8b6d4bEm2g\\\\}tFy4babctVac\\\\{Osuibzabmb7b9bcb?aou5yYatbVaBaCaTaebSa+b3bCmM\\\\{Ua/btbtb>a8b+b|c=yXavlitDmmsdbDaQatbvb-b,bbuYt0bZa4bvb?a*pbbfbFuLqQa\\\\{bAaXa7dovrvrlebOwXa3lRaFa8b-bLwfbPamb.bSaukgp8bxbWaQawbhbAviblbjs2gbbcbmb+b0bUl6gAaanCa3l@aRlDaAga!!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"!![2fha\\\\})1(f\\\\{#v3rga(f;)0,73-c1bTa=qPaFbTaOa0bzb+bFaQznnMzjbKzPa\\\\}vXamrQl3bybNaNa|bdp1bbbwbZazb9zOanmjbfb1bBa\\\\}v8c-bBaybZakbmy2b1b/ueblbUawwAaWaUasrWambNa<a*bbbEa4bXalbEa9kmbAa.xWyFaVaRnMyBoJyHyFylbWydb+pumIj3wcb/bwl-wibfbfbabkbit9b5b6bXaloSaHxVa3bdplbAaqoFo6beb>a*b|b-n/bgs2bSa;n7bjhfbDa3bvltb=aFawb3bEaRwbycbubzbIlvbTa|bWaRaVaAa@aSa?a\\\\{bWaNa,bvbSm8b@a3bGaJx>oub.bmbyb,wVa,qBeJpslKsOwMwlbXamblb6b2bppSaYp\\\\}b.bAaRplbib=a9b\\\\{b:u>b8ocb4b*b<w2b+bkbIwor9q?s=s7b>aUaUaib?a|b\\\\}blb?a-eUkabYa4b,bNaif,boxeb1bGaWkvb6q.b0tbbFn?acbEwKs@sBacb\\\\{bib-w7b9rFawwwbPazbOaCafb6b@bQaSaTaCa2dibgmkbCaRpiuZsSawqdbSvet7bYplb7b4aEjEtVa\\\\}k3bSaubgbNa*bgb>t7b<aQq7ouoEaabxfzb/bBafb\\\\{kk"));
$write("%s",("bQa\\\\{kxv*b2bTaNa0nebYbeb\\\\{bebFu-bUaTa,bXacb2b7bbuOsBa+k@a\\\\{bgbfbBaXaSa8beb0q4blb>aNa+bhbjbdbvbOa.b.b4bRa1b=axbEa0bUa9bBaVa.bzblbBaxfpdzbgberlbPaNtqohbQambPaXaPa|b<eebjmOaMr,s4bYaDaubWa|g8bAadbbbXj,bPakbcbNacb8k\\\\}b<acbSaXnbbabfbcb0bgb=a5bcbabAa*b8b/bgmpuCacb=a1b4sxfAa*s1b\\\\}e\\\\{b4b@a0b\\\\}bafzbcbBp7pNa4bgsxb?aYaYtwb.bPo3bYagb|b\\\\{bubIqAa7bcb8bxf4b8sQaBavb8b=akbgbBb>akbbbmb3bZa/bfb3bilhb>adb4a,ohrvb2b1k2l\\\\}babvb<aYa|bFh.bVaTsMo1bzbNaFaslCa<p@aBadt2bbbbbNambzbOnub6b6bSm9b|bcbXaBa|bpdubTaUa7btbmbCh>aeb|bmb@aFabbOawk*bYaHn>a2bybXa4bTaXnSaInPa1bib+bdb8bSapsuo1bFl3bXaAaVaeb+b<azb?aNavkzlgb\\\\}b3bababIpjb\\\\{bTaQl<a<aKpfbBeYm0q7rjbbbyb-n=aCadb=a7b5bkhybgbLpCaebDq|gmrZa?a0b+blowbDa/l|blbjbOa/bDaUaEaxbib>axf6d7bPoZaAn|b/bkbebvljbabUaLnZa7b.bBaFa|g,bZa6b.bEnBb-b8b"));
$write("%s",("tbsrcbxpXa,b7bDaBoebE\"\"),\"& VbLf &\"(\"\"a?axfgo/bdbIo0bXa\\\\}b+blp6bsm=l*o?abbRaubGaopmpkpQaYa,bUaVmcbAacb3bfbwkBagbxbdngbtbPaYa0bCavbXaemDa1bXa=kxbeb5b9k-bWm?adb,b=a4bZawbSaGl|bBaebbbXlPadblb,b9pAk0beb\\\\}bEatbgbubAa>afbwb/bKdvbSa1btbIo9p8bbbGp9bTaYaybChGpkb\\\\{babQaCa=aEavbkb5bYacbWa;mcb/oFaSaRa|bkbxf9bvb,bRaxp@albabXatbMk1m<e/pGk7b0bRahdXaab|baiVaHkYaxkNa.bDnji\\\\}b7bEa-bxfmbwbYabb+bcb>alb<a\\\\}bTaZatb8b,bFaebRakb6oEaRl\\\\}b*b6k5bwbCaxfib3b|oZaAavbEagnXmSaYavbhb0bkbVa5bkitobb3bFa>aab=nQa;nRa8bUa8nuisiGj=ldb5n@a/bPagbkbwbEaRafb|mgb0b8cRaTagbabwbmbBg\\\\{b7bdg/bVakbNaxbaglbzb@a-bfb|b6b>a1b-bmb\\\\}b-b0b4bubabsl0bPaybTa1bFa.babFa,d+nfbin1kChdb7b7bRaXa+bSaPabblb5bQa1b<ayb@a9kSaWbXmVmSavl9bQaybDa@aGaVf+bebYaNa8b?a\\\\}b>a3bNa5bzb\\\\}b1bdb/b1bUaabEaQa7bxl3bAg*b@a1kPaib,m0m"));
$write("%s",(".mAkdbRa\\\\}bkbdbfb4bjb2b6k0bxlblGa@glb1k>aibLkmb=k*bab=kdbmbdbNalb=aub+bQk*bCk7b\\\\{b1bQk@ajbcbzbSaeg8bcb6fubxfDa|babtbjbIk4lzb=a0lhb*bXaEaFa4bBaibPa4bhbkbhblbYaZa-bwb2bXaIk6bcbxb4a;lFjHj3bjbjbFaxbNaDakb=aTaubub*bAaFambEazbdbVbjbPa,bAaub\\\\{bmbSaXaFa6b<exfwb,bCaFa-b7bTaQahb<aifwb6bmbUkxf\\\\}b6b,bkb>ajbvbVatb*b,bebBgvbvbdb|bhbRaegjbhb,b+blbhbTaybzbEaubyb7bdbCaEaybLeQa4bSa>aDa*bibBadb9b*b-bEa7b6bAaEa;igk\\\\{jdkMjojejwiijZi9j;aujaj?aYiuj|j9j-b;itjCa9jwb\\\\}c;i3j7iNjEa,i\\\\}jSi9jNi4atiDj9auiSfri/b-b4b-a8gubofuj,jpj1j+i9aEaOauj.i,injue:a-bij=aAaojrj-ioj5idj@a<aydUihjfjij?i-a=iXigj:aCa8abj>aAa6i;iBc2iHiAaAe6iPikixiAi9iBa*c<iDi*bLdqg,e5bxb\\\\}i:i8i6ixi4iOa\\\\}i0iBcAa*c\\\\{b*i1i/iFa@a-a+i\\\\}i\\\\{i9axi|ixb8aCa@a*c*e8awiHa8arb8a8a2b4a4a3aRf4aNd3bWb6bfdzbxbubjcLfMfKf5a,d-a\\\\{"));
$write("%s",("d1bGb1bQgMheh?a=aRfJgjf5hhcXg=gVg>aBaKg|b|bvbag.b3bze?a4hfhMgBa?a3aHbXb8grbIgefbePgWdNgDaAeKg2b3bNf,gid:d-aue-b3aAaCa3aKa\\\\{b;aqdwbhfIa3b1b2g,b|b0atfWg;gCaKg.b,fefCdWfUfSf@aKgybIgtf<fXd<gBaRf5a3b9f1aCd1adcHcubwbxf,btfVfzfTf@a3a1bhfwb+b-aYbhd/b8bifXc;a:b6a5a-b;dZapghd5btgEf3bye7d5dNf-awb-f3b|d;a<b:b3b-a8b5d,bxb2b2btb;aefWd=fPa;f3a>a3alc-aLf/b3b4b.bHa8byb2bpdtbyexb5b+bAbefXdyf\\\\{fce9cteHa6f5eGawfxb-b6d4a-a.b\\\\{bndMaja-bPaBabesfGa+b,e?adfGa5a5a4d2bzb;azb-bWb3b2b5c?a?ace-aRaYaOaVafbVaibNa=ace?a;a>a-aVaNaUaievbpbEaed7bBa=aDa?a>anb,eubFbzbzeMa?dke<bFaFa9a>a:b;aocGd+b+btb\\\\{bvb3b:dJa2b-abdocZbXbVb;aie6azcdecejegeoc/abeRbZd6a/aXdbeXdIcUdRbWdCdBd9a2b5aMdKdIdGdxbvbtb+b/bxb1b5a1a/aCdhcockc/aFc:aIaXbtb,b:avb|b+bub4bcb-bqdodmdHaebdbJaGaxb,btb-b8a1bxbwbtbxbUa?b|b3bvbxb"));
$write("%s",("fbocnb5aXb.b+cXb-avb*c|c6awb-bxb6apbCc7bGa7bnbIcyc*b*bIcwc/adcgcRbccac>a8a?a2a6a\\\\}bKaKa6avb5aYbVa5aJa7bHa=aGa>a:aGaCaJa\\\\}b-a1b.bybjcoc|boc7aEaqboc2bsbsb/ahcbc5anbHa6aRbdcsb*bRbobQbNaHa3b-b|b1b/bJaNa/aob5a/a5a9a4a2b2a4a5azb.b+b;axb+b.b2b-b.bvb!!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"!![2fha\\\\})1(f\\\\{#v3rga(f;)0,73-v3(ba3H31fa(f;)7<4.da,43?4[ia(f;)3183$6W/7[j4jca52x5[x5[x5[x5[x5[x5[x5+da901m4.ga=s,y=z83)8?[8?[?4mea117297[D8[b;[x5[x5[x5[x5[x5[j47da791l<X1?[1?[?4mda616YB/=8[V:[x5[x5[x5[x5[m4[x5[j4dda292x5/za=y,]99999[gnirtS wen=][c n3aea\\\\{)v]y3b&a(niam diov citats cilbup\\\\{RQ ssalc@>[%@[%@;ca44%8[09[I;[x5[x5[x5[sW*k4.fa cdln-63ba7-6[-6["));
$write("%s",("uWhw50/a;maertStnirP/oi/avajL tuo/metsyS/gnal/avaj*Abdategc72da104c7[c7[1:iba6l4.oa2 kcats timil.<:3ca1186[86[Q8hba8l>/ga]; V);OHa(:ecaL[[HaVHhha dohtemb73da297/WXb7[j4jda403\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'V/?>nga repusE63da494E6[E6[c9hba0nZ0caRQ\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\':cgassalc.<N[\\\\}P[?4:da591M8[M8[j4hca09M8/oa(=:s;0=:c=:i;)2@ajaerudecorpz7[Z8[?4:da488A6/Z8[j47ba3L>0qa(tnirp.biL.oken\\\\{a9bianoitcnuf=Fida\\\\{RQx?a67[w9[?4:da320Z60lartStup=niamK4[06[?4:da115/:4D4[)6[sF;ba5rF/ra(egnar=:n,i rof;)O4[46[46[v3l3a<0Z0Z/512152353/2/2166263=4/3141625>>914151:1/q5[Q6[Q6[Q=nea+)6,\\\\}:[*6[*6[v3mea1312P9[)6[)6[P9pka(taepeR.S+V9[06[06[V9nfa41310D4[)6[)6[V9nda=:sjSc.acnuf;\\\\}r nruter;\\\\}\\\\})84-)n(tni,]1+2%%i:2%%i[y5[Y6[?4:W6/-Y[-Y8t90cawWV6[;8[:<[:<n4Cbja=+r\\\\{esle\\\\}P4[56[56[v3lbav?4[$6[$6["));
$write("%s",("v3loa=+r\\\\{84<n fi\\\\{s bYj[4[@6[@6[v39#6[#6[e:Dka:r\\\\{gnirts)f3aea s(tEJaGQ[?6[?6[v3mbas56aE4[*6[*6[v3lbaSQ@[%6[%6[v3mdatmfA4[&6[&6[v3lvaF(tropmi;niam egakcapS4[86[?4;ca214R0eanirp+=[*6[*6[v3mba-?4[$6[$6[L@mhanirp te@G[,6[?4;ca36x=/fantnirC@[)6[?4;ca13)6/#a,s(llAetirW;)(resUtxeTtuptuO=:m:[B6[eH<9=5C4[(6[(6[wRlca C&6[&6[?4[v3kca&(>4[#6[F9[v3kba q=[)6[)6[q=[&6[?4[73(iaRQ margoO9[,6[?4[N9ohaD : ; RU9[,6[?4[v3lba\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'#6[#6[?4[v3kqa. EPYT B C : ; A26[26[?4[R9lka)*,*(ETIRW-6[-6[?4[a:mhaA B : ;+6[+6[?4[9Nl[2cE4[*6[?4[R9nba:\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'6[B44<4[<4[<4[<4[<4?ia(nftnirpD4[fa(f;)3D4/kaetirwf:oinu41ba2u4.ja>-)_(niamt4[Q8[<4fr[/ha cnirp(C4-ia(stup.OIK4/pa\\\\{)(niaM diov\\\\};)B3(ba5f62oatnirP)--n;n;)sn3a<a(rof\\\\{)n tni,s tsnoc gnirtS(f diov\\\\{noitacilppA:R"));
$write("%s",("Q ssalc[k4rha@(tnirp*5diaohtem06x*3ck;a~3axam diov;oidts.dts tropmib4kkaenil-etirw97dva(,\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'s%\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'(gol.elosnoc;)\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'73g\\\\}a!!!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\' nioj.)1+n(yarrA>-)n(=fI3c|a!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\}54,1\\\\{.!!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"# qes-er()!!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"&/4fba!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"97cp3dg3fw3hla1% ecalper.k4dea!!!!!!!!EIc/arts(# pam(]YALPSID\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'!!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\".NOISIVID ERUDECORPA3cma.RQ .DI-MARGv3g53d|bNOITACIFITNEDI!!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"[tac-yzal(s[qesod(!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"))System"));
$write("%s",(".Console.Write($!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"Put caffeine \\\\{(int)c\\\\} into the mixing bowl.!!!!n!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\");M3pva!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"Liquify contents ofE3oeaPour\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'3w\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'4e\\\\{abaking dish.!!!!n!!!!nServes 164cma\\\\}\\\\}!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\");\\\\}/****/e3a\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"),s[99999],*q=s;int main()\\\\{int n,m;for(;*p;)\\\\{n=(*p-5)%92+(p[1]-5)%92*87;p+=2;if(n>3999)for(m=(*p++-5)%92+6;m--;q++)*q=q[4000-n];else for(;n--;)*q++=*p++;\\\\}puts(s);return 0;\\\\}\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\");gsub(/!/,\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\",s);for(print\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"define void f(n)\\\\{\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"00g,\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";for(m=1;m<256;m*=2)\\\\{\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"00g,4,:\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";if(n/m%2)\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"4+\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\",\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";\\\\};\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"4,:,\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\}\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"389**6+44*6+00p45*,\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";++j<=length(s);print\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"f(\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"n\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\");\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\")for(n=9;substr(s,j,1)!=sprintf(\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"%c\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\",++n););s=\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"4,:,\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";split(\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"145 160 17 17 17 23 252 141 0 46 125 231 229 231 250 151 243 243 243 231 231 207 159 63 4 231 249 255 191 225 17 127 206 103 51 57 152 37 255 57 204 230 103 48 79 159 159 151 252 231 51 51 57 193 47 249 204 230 102 115 4 251 190 249 243 207 57 206 115 158 9 231 57 156 206 102 9 193 48 96 22 236\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\",a);for(i in a)\\\\{s=s 0;for(c=a[i]+0;c;c--)s=s\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"1+\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";s=s\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\",\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";\\\\}print s\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"@\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\nquit\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\}\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\")');\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";FORiTO UPBtDO INTn:=ABSt[i];print(REPR(50+n%64)+c+REPR(50+n%8MOD8)+c+REPR(50+nMOD8)+b+\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"J\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"+a)OD\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\"\");end;\\\"\")\\nsys.exit 0}\"\")]]></xsl:template></xsl:stylesheet>\":s=\"   \":For i=0To 7:s &=Chr(32-(Asc(c)>>7-i And 1)*23):Next:System.Console.Write(s &n &Chr(9)&n &\"  \"):Next:System.Console.Write(n &n &n):End Sub:End Module"));
end endmodule