module QR;initial begin $write("%s",("let s=(\"Module QR\\n\")\nput=s\nprint\nlet s=(\"Sub Main()\\n\")\nput=s\nprint\nlet s=(\"Dim c,n:Dim s As Object=System.Console.OpenStandardOutput():Dim t()As Short={26,34,86,127,148,158,200}:For Each d in\\\"BasmCBBBCRE`F<<<<C<`C<B`BBD#CXwasi_snapshot_preview1Jfd_writeBBEEDCDGECB@IUDHmemoryDBH_startBDL|DRBAC BAJlACA4RB9MiCD<AERCA>D!BE@ABRCABRCABRCAJ!CE@ B-BB CACk:CvACqRC COBMADRCACRCADRCABRCABRC BACj:B-BBOBMADRCADRCADRCAFRCMM}CBABM~(BBBCBBB,BBBDBBB0BBBDBBB4BBB=BBB?BBB;BBB ...\\\\t..\\\\n..(module(import :wasi_snapshot_preview1: :fd_write: (func(param i32 i32 i32 i32)(result i32)))(memory(export :memory:)(data :\\\\08\\\\00\\\\00\\\\00$:))(func(export :_start:)i32.const 1 i32.const 0 i32.const 1 i32.const 0 call 0 drop))\\\":c=Asc(d):If c=36:For c=0To 11:s.WriteByte(If(c Mod 3,Asc(6"));
$write("%s",("43811.ToString(\\\"x8\\\")(1Xor 7-c*2\\\\3)),92)):Next:Else:n=(c>124)*(8*c-41532):Do While n>127:s.WriteByte(128+(127And n)):n\\\\=128:Loop:s.WriteByte(If(c<125,If((c-1)\\\\7-8,c+66*(c>65And c<91),t(c-57)),n)):End If:Next:For Each c in\\\"<?xml version='1.0'?><?xml-stylesheet type='text/xsl'href='QR.xslt'?><xsl:stylesheet version='1.0' xmlns:xsl='http://www.w3.org/1999/XSL/Transform'><xsl:output method='text'/><xsl:template match='/'><![CDATA[sub f(s$,n)print(s$);:for i=1to n print(\\\"\\\"\\\\\\\\\\\"\\\");:next:end sub:f(\\\"\\\"write,format=\\\\\\\"\\\"%s%s%s%s\\\\\\\"\\\",\\\\n(\\\\\\\"\\\"\\\"\\\",2):f(\\\"\\\"write{-}{txt}{echo -E $'(\\\"\\\",1):f(\\\"\\\"\\\\\\\"\\\"with Ada.Text_Io;procedure qr is begin Ada.Text_Io.Put(\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans B(Buffer)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f("));
$write("%s",("\\\"\\\"\\\\\\\"\\\"trans O(n)\\\"\\\",2):f(\\\"\\\"{\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"B:add(Byte(+ 128 n))\\\"\\\",2):f(\\\"\\\"}\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans f(v n)\\\"\\\",2):f(\\\"\\\"{\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"O(+(/ n 64)107)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"O(n:mod 64)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"O v\\\"\\\",2):f(\\\"\\\"}\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans D(n)\\\"\\\",2):f(\\\"\\\"{if(< n 4)\\\"\\\",2):f(\\\"\\\"{f(+(* 6 n)9)48\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{if(n:odd-p)\\\"\\\",2):f(\\\"\\\"{D(- n 3)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9"));
$write("%s",("):f(\\\"\\\"\\\\\\\"\\\"f 27 48\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 36 11\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{D(/ n 2)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 21 48\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 48 20\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans S(Buffer\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"STRINGz:=REPR226+REPR153,a:=z+REPR166,b:=a+\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"2\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"+z+REPR160,c:=b+\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"8\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"+z+REPR165,t:=\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"class QR\\\"\\\",2"));
$write("%s",("):f(\\\"\\\"{public static void main(String[]a)\\\"\\\",2):f(\\\"\\\"{a=(\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"write(\\\"\\\",4):f(\\\"\\\"'implement main0()=print(^1^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"BEGIN\\\"\\\",2):f(\\\"\\\"{print(^3^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"echo ^1^\\\"\\\",4):f(\\\"\\\"'f(s)\\\"\\\",2):f(\\\"\\\"{System.out.print(s);\\\"\\\",2):f(\\\"\\\"}s=^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"389**6+44*6+00p45*,^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";for(c:(^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"#include<stdio.h>^8^"));
$write("%s",("nchar*p=(^15^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"Ra#include<iostream>^16^nint main()\\\"\\\",2):f(\\\"\\\"{std::cout<<(^31^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"class Program\\\"\\\",2):f(\\\"\\\"{public static void M83abbSystem.Console.Write(^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"Quine Relay Coffee.^64^n^64^nIngredients.^64^n^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");for(int i=9;i++<126;)[3pva$^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",2):f(\\\"\\\"{i\\\"\\\",2):f(\\\"\\\"} g caffeine \\\"\\\",2):f(\\\"\\\"{i\\\"\\\",2):f(\\\"\\\"}I3b54rja^64^nMethodv4f#aeach(char c in(^6"));
$write("%s",("3^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")))^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^32^[2al3dp3c[2cs3c,3l[2k@3kqa^31^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")s rts(ecalper.h3eja^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"     53c4a SUTATS(egassem^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"rts(nltnirp(])]^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\".NUR POTSu4cba.C3dh3dX3bba[65bX4df5lp3lna\\\"\\\",2):f(\\\"\\\"})1(f\\\"\\\",2"));
$write("%s",("):f(\\\"\\\"{#\\\"\\\",2):f(\\\"\\\"};)06xt3dba;+3nna3(f\\\"\\\",2):f(\\\"\\\"{#qp]^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'[p]#3sv3r23)ga7(f\\\"\\\",2):f(\\\"\\\"{#.33)ca51h4-ba1S4w23F?7d33&r7u53sda,4353.ma^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\"));
$write("%s",("\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"' D ; EYB RCL4/v4+ja36(f\\\"\\\",2):f(\\\"\\\"{#DNEm4[m4ada. A~5[p4deaPOTSn4[#5e~5[o4boaRQ margorp dnex4[x4abaS*5[m4c2<[ca91j4[j4eba&%6[l4bgaS POOL)<[:7dba^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'j4[j4[j4gda&,)(6[?>cga. TNUO<7[s4bfa(rahcg:[(5dgaB OD 0B>[t4cca&,,<[,<aca)A36[;=e6=[.6cqaEUNITNOC      01z4[c9c,5[W8dK7[aGeeaRC .p4[p4aka,1=I 01 ODt4[TKecaPUq4[/I[6<hva;TIUQ;)s(maertSesolC;^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\"));
$write("%s",("\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'Ye%4Rra744(f\\\"\\\",2):f(\\\"\\\"{#tiuqn\\\"\\\",2):f(\\\"\\\"})215>5[qa^32^\\\"\\\",2):f(\\\"\\\"})959(f\\\"\\\",2):f(\\\"\\\"{#n\\\"\\\",2):f(\\\"\\\"})420pY4d8,ba8AAbg8[da304zY[O7bda218lK[wL[j4ldamif+6[ga)91361\\\"\\\",2):f(\\\"\\\"}5[,6[j4lbat(6[(6c%a315133A71/129@31916G21661421553/04[04cva%%%%\\\"\\\",2):f(\\\"\\\"}*+1%%%%811 -\\\"\\\",2):f(\\\"\\\"})48\\\"\\\",2):f(\\\"\\\"{3bhaj:+1 j@34[34cbawm4[m4cl4[l4cbaWm4[m4cba\\\"\\\",2):f(\\\"\\\"{m4[m4cva)(esolc.z;)][etyb sa)t=[#>[j4[<6hea3289m4[x5[j4lba,l4[w5[j4hla!\\\"\\\",2):f(\\\"\\\"})46(f\\\"\\\",2):f(\\\"\\\"{#~~v4[%5[j4hea(rt.o4[z5[j4hba)A7dda\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"};l3efa~~dneo3hra~~~~PUEVIGESAELPnr3ala~~1,TUODAERw3a63j$a(etirw;\\\"\\\",2):f(\\\"\\\"};u=:c;))652%%%%)u-c((||13jda#-<q3jda||i)3mhaBUS1,ODs4qka)3/4%%%%i(N4cx5kU4xPa2=:/t"));
$write("%s",(";2%%%%t+2*u=:u\\\"\\\",2):f(\\\"\\\"{od7 ot0 yreve;i-=:u;1=:+i\\\"\\\",2):f(\\\"\\\"{od))1(evom(dro=:t elihw?s;)s*45oi5vv3jd7dladohtem dne.s3dganrutern3d~aV);gnirtS/gnal/avajL(nltnirp/rZa|atnirP/oi/avaj lautrivekovniJ3d.4j[2cib\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"};0=q;)]q[c=z(tnirp.tuo.metsyS;)0(tArahc.y+z=]++n[c;y:]q[c?n<q=y\\\"\\\",2):f(\\\"\\\"{)0>2%%%%++i(fi;48%%%%)31-)i>3c&as(+87*q=q\\\"\\\",2):f(\\\"\\\"{);47522<i;(rof;n)rahc(+K4r[2k*3&oa=]n[c);621<n++r4aqa0=q,0=n,0=i tni;N3&kc1m4asdRbQehmxfvfamRf<bedPdck\\\"\\\",2):f(\\\"\\\"}b;agb-a|dzdxdRfGb8aqeRdYd5a\\\"\\\",2):f(\\\"\\\"{b2bGi;agb-epb>a8adewj>aJaRaAdteFbaeIfOa5aac2gJY6f9a<+4aLa7a;a4a<aPhnnkdxd;aNa?c6a|eebHaFaIaebzeJaeb9a/a6a2dQbUe-f2a-f9a<+5d6cRbC3g7c-f/aof0fRf6q7esko62e6aRa;dNaxbogI+Gh;aTapc4aLcEeyiof6amc<byg-fFmsbvh\\"));
$write("%s",("\"\\\",2):f(\\\"\\\"{2WfybxcxcB@UeAa2a6a\\\"\\\",2):f(\\\"\\\"}g7a6a@a\\\"\\\",2):f(\\\"\\\"{g:a?aMbKaKa6a?e:a@aEa2a|gZfMbbgli>a:b1a-glnUf\\\"\\\",2):f(\\\"\\\"{bHa4atcEi<7wbJ;+bfkJ;\\\"\\\",2):f(\\\"\\\"}bJaMa\\\"\\\",2):f(\\\"\\\"}bJaq|Ec-bJaJaUa-bJaMdJa8b9Y;a8b/vKa8bSa,RT*ZtnF?u<79bs3a\\\"\\\",2):f(\\\"\\\"}a\\\"\\\",2):f(\\\"\\\"{8,RU<Sa,R<7wb\\\"\\\",2):f(\\\"\\\"}bJaLaJa8bU<<7j4coa8b<74b<7:bJ;+b*4aiawbZtJaHa\\\"\\\",2):f(\\\"\\\"}3a=3a-aHaJaFdqN;a8b5;:aUa:a9YviSfQfNm4ap\\\"\\\",2):f(\\\"\\\"}sbsb2be3^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'maviDa-a|b?+-aD6aua?aGaUe>a/j\\\"\\\",2):f(\\\"\\\"{gKaKa|gZf(6cgaagHkkg,6esasbvh*b-a/bxcHa|fDle3c0c\\\"\\\",2):f(\\\"\\\"}b\\\"\\\",2):f"));
$write("%s",("(\\\"\\\"{gph\\\"\\\",2):f(\\\"\\\"{gvg1a-g\\\"\\\",2):f(\\\"\\\"{bHaDlRf-e:a:a\\\"\\\",2):f(\\\"\\\"}bHa?a\\\"\\\",2):f(\\\"\\\"{gJa\\\"\\\",2):f(\\\"\\\"}b5aAdte@a1a-g0iDlxcpb7anb2b:b\\\"\\\",2):f(\\\"\\\"{g2f7k@d-aIfVkxcHalgjghgal-aUf0ixiRf-f-gSf|fDlzeSgxiHaTk;a/aDh<b+hWh<apb/aDhWhnb<ags:b\\\"\\\",2):f(\\\"\\\"{g/aDh-f-g+gFa,i|b1ali3b:b\\\"\\\",2):f(\\\"\\\"{g9hHaDlHaUe-iCe|bxc3b0a:b\\\"\\\",2):f(\\\"\\\"{gIa|bzeJa|c5b#aQbxi<b=a-aAn*c3bxdUe=a-a?aaB9ai3edb2bMa7apb3Aphnhlhjh9apbqhohmhkhKcdc/bPcgfvfOhJh7a3A.l,lMaAn*cEc,dJa>a2aIfUjMgMa?aaB<i+cbi6a/3iYaxdHQvb8g/aDh=apiRalbOaCdlbrU3-@Zpi0k6a7b5aTkRfwbXjUe2bAdwm|\\\"\\\",2):f(\\\"\\\"{-bhcloOiOihq0c/bxd;a<hJj-?aea6a2bR>e\\\"\\\",2):f(\\\"\\\"}cnCkO6a-o2a5a+knI\\\"\\\",2):f(\\\"\\\"}gEhgl/b-bOi6aUh9mHa1dmdLhRfNl7mHa:eNl7myk;almQaCORfmG<b3bxd6aIh:l5a*jUVkivftfv\\\"\\\",2):f(\\\"\\\"};a9jcc8bfbpbubldic+d,bnbpgPjNjEc,d"));
$write("%s",("0kfl6m<b<b<b=k:b3k<b<b,cBk?k7b-bBkEa<o3bDdzlMi9a7b6g-a5btx,cBk=a9a7bubxbs3e33eca:k33eea.b8fE3c33ifaJb7bd^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'3fka:k=o6q9ai8)3cmakiolKj9l,cBki3aCa-a+bhh.bfh,cBksbHa\\\"\\\",2):f(\\\"\\\"}gmkMlkgKlMk;kCaLi6a0kflXkik6a6lWlPkUlxl<bzebDc93gea1lLi+3edbF1E:VR0c4mqk2m0kfl?l=l3a6a<bki>j/yE:VRNT2a2amGVkPl0iwbXjRf@a>anc:e7b5aWf=anbVkybsl5a,bJa6a3Aa%aub9h5aUgwbXjHa:e-b9a9b9adlVkyg>am3a\\\"\\\",2):f(\\\"\\\"{a@a@aVkyg@a>a:a|b9a0b9a@a>a#Ca?a>e|bPg9bJa0bVkyg-b9adl9aCaAaJa9bVknbJa6a|b5a,bRf:e-b.lw+-a,<a&aTvE:VRvimGyg8bAdGh-amG*bD5-amGyg7s3heamG?a,6cca.jt6a5amGKc>irPxd6a-b"));
$write("%s",("9a8b9a7bJcJayb>akvki>aJa*c@dxc?bo\\\"\\\",2):f(\\\"\\\"{o3a3a-bEmteUe@a>a<a2b5aDcxbvb:atcJaub5aEcxbw2|\\\"\\\",2):f(\\\"\\\"{-bVgE;aeaJlHlS;aT:akamG7esktjpkr8g%eTlRlpb;awbXjsmmGmGd?lAjO38jnumPnuo@mUm1o/oCnEo@a;oQ,L*hczq@6\\\"\\\",2):f(\\\"\\\"{iqIkOpC;ZGW4.0GKykiO6JtjbLo3volq|Val0/,Wrlbuski8WCa+M0>Zafpk+lb=rZafpypp\\\"\\\",2):f(\\\"\\\"},bfb-bhvQa-bLoH46b1bgb<a>alhR9ZaL*UZHS>aG6JAEEF?m\\\"\\\",2):f(\\\"\\\"{2bgb=aFajb>0Paoq??DaIw@qoqm/5vLtabJu1bDa,b7b<3hbm=lbI|BaMF\\\"\\\",2):f(\\\"\\\"{bUaTJ9-abE=Ba/\\\"\\\",2):f(\\\"\\\"{RSoj3bEp,bZMR9.rabh8HY69Zqo1h*WIjbP2fKub/b=a69-2q7\\\"\\\",2):f(\\\"\\\"{bq|UDDrlbSHWsybNSfbyyYz5YY9C+3bFs5zwSh3|bcblP5b-Djpjd<@9jmb|b7bDBwxUa/>>6e$d+.*b<aYaW\\\"\\\",2):f(\\\"\\\"}jB>;wSoG4qIz@6g7U\\\"\\\",2):f(\\\"\\\"{2*i9=xp.lb\\\"\\\",2):f(\\\"\\\"{PTav.>ippcmuwki<<1z6.3-|sK0EyrgT<dv-b5pFiFUZa\\\"\\\",2):f(\\\"\\\"{bXzCplrCtJ"));
$write("%s",("wB7Ayjb1,6CcykiQC9Gz.+po.ScNaJv4.G8SaD?8rR|5/N5+4LXZbD?.\\\"\\\",2):f(\\\"\\\"{r\\\"\\\",2):f(\\\"\\\"}ywo\\\"\\\",2):f(\\\"\\\"{vtZA|bwLYafCCa.E7bD?<GI9T4Y:lboA8\\\"\\\",2):f(\\\"\\\"}lYSw3wSw2bnp9q7;EaWa4PJpf3@azs6uYpmb5Y\\\"\\\",2):f(\\\"\\\"};9zXaybzbHrPO/bZamb|;NFbpFB\\\"\\\",2):f(\\\"\\\"{bg5?xqyebaboAFA9bEa6uZo5b9+cp>sEa,6e~d5b>v*t<a,bdu6bP>Cp0Mn+3*2byLCVAVFr\\\"\\\",2):f(\\\"\\\"}r@s1VB.t8Ru7\\\"\\\",2):f(\\\"\\\"{2z?pNU:RH2?phbWrFZ1PzbX>zB@aFUlYIXbXxqSaQ2Lo@=-<Da55y.er>ai/Saop;sCaQo/b0bo8@W1xkh,5B</rBIouhb?aEZztkijzepgp*bjbYD1/krEa>aa82*?U,\\\"\\\",2):f(\\\"\\\"}Da<U@aTaer>agRHuo8q*o*q;/vL\\\"\\\",2):f(\\\"\\\"{/v;w-1jb?nkNEpDaN-Ca?L=a-bkNy|UCVa/,lb>Agp2bdUVadpmbwqEacb+.3AAwNacb+.q3exNaZ74;\\\"\\\",2):f(\\\"\\\"{btx*6e$bZaZuPQiFiuwqEa51J|wb5pW:B.Q2=T+sB.;wopbHZo\\\"\\\",2):f(\\\"\\\"}bZLEaSj-1tGw:?x<p6bm*Ea\\\"\\\",2):f(\\\"\\\"{bdbZoo7\\\"\\\",2):f(\\\""));
$write("%s",("\\\"}V\\\"\\\",2):f(\\\"\\\"{bwqEaE||ufpkbfbZuLX3vIzZu9b9C=G?xQ;prFF\\\"\\\",2):f(\\\"\\\"{3s5aLb4\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{3ubDa8;Zo5bX>J8RDEa5bX>VrHyGDubVr+;gbCaL:IS?a;3Ea4q5bDSC>TadyylJ8<aGq:SgbVXsIXoh.U\\\"\\\",2):f(\\\"\\\"}tshbowDacN:>Kyub,p/b25=atKg>hbt9/p-phbf3c4TlX>r1qS0l0bwSLq1lW5dx9+=aGqXM~6eoatbc4Tl9+<aPR?x+3cMcDaH<r.hbWyG>fJ3H3+hbRatb>ahbTl/p-p-H?Reb0pb20XqS+-3Oi>qqZaFa|qEaSzeQUp5bsq2,+r;zh8j6D6/rSZ.r6j0>7qKtDrlb>=6|Cq<W,R>I<Ifx*qK\\\"\\\",2):f(\\\"\\\"{5tswGtsw|bhbmbFv>5+babL0=aTF@a@amsK36zAnl7hb-qlbk2Sahb|yj:Oa6wab?e?C1Bhb2X<71Bhblb/,8\\\"\\\",2):f(\\\"\\\"}A0.41CCLh.Sl=LK/TaCx2I4PguMpWazztc@1$4ciaub+|zbA|$6ewaksz:x:6.yb+bBa:vzbW\\\"\\\",2):f(\\\"\\\"}bKi3qPc5bq8W\\\"\\\",2):f(\\\"\\\"}bKi.vb=x6/\\\"\\\",2):f(\\\"\\\"{GRC3xv\\\"\\\",2):f(\\\"\\\"{Ear\\\"\\\",2):f(\\\"\\\"{3=B2ONMpwb6+MSxsDrNU:sDa.b.bWIWr\\\"\\\",2):f(\\\"\\"));
$write("%s",("\"{OY9zthbubhpr|kpB\\\"\\\",2):f(\\\"\\\"{xhl15V@aHr4tGpm5jbNaxbDal;vb8b>=h\\\"\\\",2):f(\\\"\\\"}tb|wqx=<UFTaib>3*Yf3Gu+q6W|\\\"\\\",2):f(\\\"\\\"}gsd|Fapu=6Ixcr0bG+x-+MFB,Rf\\\"\\\",2):f(\\\"\\\"{1b7bbjebh1ibYaSaI\\\"\\\",2):f(\\\"\\\"}KtOaH\\\"\\\",2):f(\\\"\\\"{Xaj\\\"\\\",2):f(\\\"\\\"}E6-qRI@U>UbyTWQt\\\"\\\",2):f(\\\"\\\"{yubzbRok/PaGYfb3w2,ic\\\"\\\",2):f(\\\"\\\"}rD?5Cmb|O0-*>N>@fGg9:=sxY9babA\\\"\\\",2):f(\\\"\\\"}E0hb\\\"\\\",2):f(\\\"\\\"}bQwq?Gu;B6bubO8nyS|CaT9*:og+HZaE=hZa*v|6El0dp8;qV0boV=zvp\\\"\\\",2):f(\\\"\\\"{ylbj\\\"\\\",2):f(\\\"\\\"}ubE=GaC/x2uAhN|-6bZL7baMM:k>IzB+J-m*Gu;Bd1lbp?ptx7*b<x<:9L2bVomrZaRagbvxvb8bPt.bNaL+Muk>NysrZrM/b,+bjbR1+4ab266\\\"\\\",2):f(\\\"\\\"{SacxPXy\\\"\\\",2):f(\\\"\\\"}4qdbgbA\\\"\\\",2):f(\\\"\\\"}2btWh\\\"\\\",2):f(\\\"\\\"}UakbNVFkoutb51Swmrow><yv7x5x4:;q6>,ua/>=?a|-YKb\\\"\\\",2):f(\\\"\\\"{.t3wps\\\"\\\",2):f(\\\"\\\"{Fs\\\"\\\",2):f(\\\"\\\"{WiIuJ4dFj|g4CXPTXR"));
$write("%s",("E:VRgA+.9f-b?\\\"\\\",2):f(\\\"\\\"{,bbb1bCawbP5\\\"\\\",2):f(\\\"\\\"{b7|MYQacvUy9b6b\\\"\\\",2):f(\\\"\\\"}bmQub>a/4Ky8>3b6>,uGE>,ybAwKz1wJvB0yb-l/bBLITrS5.7bl8F9.4qy,?0b=aScnyaM=sIQPt3BCa0RztHr=WPOK*3Bublpo01u>+d\\\"\\\",2):f(\\\"\\\"{/@EvnyI:l0QaZa=z.bmQt-jR@s:r=+Muj9Ny:sz,t+wW*>f97\\\"\\\",2):f(\\\"\\\"{0\\\"\\\",2):f(\\\"\\\"}@aRxPa@abxS=9Yyb<DGa\\\"\\\",2):f(\\\"\\\"}TPW?a+bNyCtVa3w.b2X=+lb6+@+3IQaBy<KQqpqw*,,4ZTaq.R11x6b8\\\"\\\",2):f(\\\"\\\"{Xaki@\\\\\\\"\\\"),\\\\n(\\\\\\\"\\\"+ZaylopX\\\"\\\",2):f(\\\"\\\"}9G3B#=f>curKMsZabxW*jb08Val0CCyr2.D?nSHsnSD?utIU4p/@twrwTWQarS3bkd6sC7O1T45R:I6tRQU9=rRoUq+zlyjbO:\\\"\\\",2):f(\\\"\\\"}VZ-JARa;HwbT,wpZaub+j-\\\"\\\",2):f(\\\"\\\"{yMB=vy8\\\"\\\",2):f(\\\"\\\"{Xac/+bCa1b1G1\\\"\\\",2):f(\\\"\\\"{1bcW@zHrT2>aJL6/kd6sI\\\"\\\",2):f(\\\"\\\"}Q+.5aiz,Q+.5s1H52,2,+r69S\\\"\\\",2):f(\\\"\\\"}K0=6Di+-Swl3UolbAZe8Eabb\\\"\\\",2):f(\\\"\\\"}0o3eb=,Frs\\\""));
$write("%s",("\\\",2):f(\\\"\\\"{cm@+f*8-/W5-A3a/a?|p\\\"\\\",2):f(\\\"\\\"{.\\\"\\\",2):f(\\\"\\\"{2,lb4bBaGaYWfbl08L+rAL9=324\\\"\\\",2):f(\\\"\\\"}Ea5b-z/b|6e%dXpK2Jwj9<Dm22zuVdbxUUF\\\"\\\",2):f(\\\"\\\"}Vkb5pl3+bD-3v4\\\"\\\",2):f(\\\"\\\"}n8nhYaEa\\\"\\\",2):f(\\\"\\\"{bPaVX-qNawb3rGa\\\"\\\",2):f(\\\"\\\"}TxU|bs1wb/qUS=aaycKLXHrkbyrh3;ski+W8rv,L0h1Vx3,q|<Y2+zbiItwUWow6.U2UZhbjbFa\\\"\\\",2):f(\\\"\\\"{V-b:-Nahhw\\\"\\\",2):f(\\\"\\\"}8r6*8qzbb\\\"\\\",2):f(\\\"\\\"{KB9GUap;xbNa3bNUaiU1NaxbNa=<K>7.2b6b4|XqOaY1i/6Jc3Pj?fybZa\\\"\\\",2):f(\\\"\\\"{|xbgueu3?+v5b3-Eat4?4G:O4Pyy53-0vD=y5;JMFCa6|cp@rg+m5KXUaos9b3b6t.bAx?qh+LK9f/aYs4bebnF9wa\\\"\\\",2):f(\\\"\\\"{.dNaacmw\\\"\\\",2):f(\\\"\\\"{FHWl8\\\"\\\",2):f(\\\"\\\"{bE4Ua9b+-hbdbj1^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9)"));
$write("%s",(":f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'=cEc?a>1wb9GHr15<IX6rSTBSzgbgbgb+BvbL\\\"\\\",2):f(\\\"\\\"{z,9\\\"\\\",2):f(\\\"\\\"}HjOoldLQ@ams@?L,f.nSY0XtjrebrSV.eQaicbC\\\"\\\",2):f(\\\"\\\"{|u1rmb2bhC2,0:V9Mho1VtV6e7c7IEo\\\"\\\",2):f(\\\"\\\"}ZjjvXQr.@S=kKozqwvG34b<aupRX*Do0RVoqBaIEYa1uC\\\"\\\",2):f(\\\"\\\"}08vb@89Aabvx=Lzxl1kRT-C\\\"\\\",2):f(\\\"\\\"{>a\\\"\\\",2):f(\\\"\\\"}z+bwb:XO2e7c7r7Fa<WHYQ,i.1xlpPaG,tsg5,b+bwbibqvIHwvTaw=(6e5a/vwLFaLJ\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}O94bib9zXzuqFaWI?ak=d0cb@iEan9hbjb<BDCy3c<c/b@auKLh0\\\"\\\",2):f(\\\"\\\"}Va:Daz,bWAH2i*Q=cbd7l0vbRpRQZ+mji.BMw\\\"\\\",2):f(\\\"\\\"{7PF<4;Ay;,Sa@ah7w=Wa|C9\\\"\\\",2):f(\\\"\\\"}h\\\"\\\",2):f(\\\"\\\"}0bwtf1L2ab@a+bFBOU3BAagX+rTs1:\\\"\\\",2):f(\\\"\\\"}u.:xuy,w+og5Y.5+r37Vaf>e|8t9Aab6.2bxRc5hbTQHj/.BT=aJ0eU|HUums=aZBibPFNaC+s+9bCaIUywRSC+TagTV"));
$write("%s",("so*hbr\\\"\\\",2):f(\\\"\\\"}*Djx86-?yw\\\"\\\",2):f(\\\"\\\"{|k8IzR;P;0brr=1Gfpdeb?I=I8t6bGB2*<ko>fudubu5*<kNYTt@iWa3rX@kiiXvbN,T<5R6b36i*ku7R,Rf\\\"\\\",2):f(\\\"\\\"{:jAp6CKz/bA@PxDPo.cLIBAQ956C2pzb\\\"\\\",2):f(\\\"\\\"}@Pa9rt?z:U+kzIWkiGV4p=9=<;|8q6b.wwD\\\"\\\",2):f(\\\"\\\"}Q0bbbubFakL6bPw@5Pz6\\\"\\\",2):f(\\\"\\\"{y7sro\\\"\\\",2):f(\\\"\\\"{LKIULKUaGAO\\\"\\\",2):f(\\\"\\\"}Pa@4m3WIzsPs5s-JKz:wwbWa\\\"\\\",2):f(\\\"\\\"{rkbaiWAR6OC6bN56b0Ab2=\\\"\\\",2):f(\\\"\\\"}K2vxwb=k|D<IDTCaH/|bXALrlb0zIoUa|b:\\\"\\\",2):f(\\\"\\\"{1xzYrUohq/M?dyw=3rx6e5aQ20zAs2|.blbQs*bUq|bzYZh4+s*YvEZ6b6bg\\\"\\\",2):f(\\\"\\\"{>sBMzY;,*1u3eOaRa\\\"\\\",2):f(\\\"\\\"{b-0Ua4b9qo4oy4UYa@abbeu,bf9PzR|RIEZPzfbXQ0bFaKxe-\\\"\\\",2):f(\\\"\\\"}bSH@S4.8*Oa8rNaAa@ar3?3aGbU.GoDT9GBaAwY+VPQ,S\\\"\\\",2):f(\\\"\\\"}T,WID>WMSUZq*D-.Qz8qEy2,kb;\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}1,b7\\\"\\\",2):f(\\\"\\\"{1RKXUzFHv"));
$write("%s",("b3w.b;vF9I+vb5M7bFai.aHEamQ5R<af5K551\\\"\\\",2):f(\\\"\\\"{b7b/,PDxPx-6+MS32\\\"\\\",2):f(\\\"\\\"{bybM5YT@tIpI@Ms1l?rDw5.WBJZ?al85bFE9f+d+4W;Sa@MVaguTa7b-bS40GvbE,xb@t,xkPUpusPX\\\"\\\",2):f(\\\"\\\"{bX.8b4.?aL*8Azb4.Ca0xnyPaRaZB+bi:dbxbex,x\\\"\\\",2):f(\\\"\\\"{b\\\"\\\",2):f(\\\"\\\"}V>r0b.xTrNa3bn?g\\\"\\\",2):f(\\\"\\\"{.bo\\\"\\\",2):f(\\\"\\\"{1,K*LKts5.fKRM8bNa.Qm3wbI@cpFG;vXVH\\\"\\\",2):f(\\\"\\\"{lrIGTa:RgBNa/?jUKtYTM+ly--ki@+wb>ac\\\"\\\",2):f(\\\"\\\"}>s;i\\\"\\\",2):f(\\\"\\\"{EUpVa\\\"\\\",2):f(\\\"\\\"{rxwWryljbq@pq5bM5LWwbjbrw?aY1hb\\\"\\\",2):f(\\\"\\\"}b0w/CEahz1b?vJhaRFM?a3O6bzqwSki/O7sbyxvgz502b3x.R@Ms+2|-bmsi*m;4t3\\\"\\\",2):f(\\\"\\\"}?hkbd5tbq|glDfSa:R2b,wNF3r777<NF?auKL>YyI@1<lb0b+>2bw2.b.bd2Oj?aeuebF9.4OSIR\\\"\\\",2):f(\\\"\\\"}V2WGvq-2P@+EHGMVai3a/cZaJ-3s@g3rU3DaQ:5.HPhbbx/bIuuN@aTaJLgBPaVi3w9LOo/bibe,twrwmr<w2bNxr6FYPX9v-Ilb1z5z1zb\\\""));
$write("%s",("\\\",2):f(\\\"\\\"}qygbxb=sStIuQa<\\\"\\\",2):f(\\\"\\\"{ubEa=-f5yb\\\"\\\",2):f(\\\"\\\"{b\\\"\\\",2):f(\\\"\\\"{|32q>gb|b0bcr\\\"\\\",2):f(\\\"\\\"{b0wYv;Jyb?eUVtJ:2l:iIfhs+I\\\"\\\",2):f(\\\"\\\"}W*0:Ba<B+b1bCx??abfxnyccUV@+hbtsybIg\\\"\\\",2):f(\\\"\\\"{wP8OA.G|bbkJ4i.1-1bd2f>fRitdOv084BbHewhb?hxzvx=,FYubfx5qE.7wGEbUw\\\"\\\",2):f(\\\"\\\"}eDIu/4JY\\\"\\\",2):f(\\\"\\\"{IXwQaD\\\"\\\",2):f(\\\"\\\"}kbY|m*0Gabms3bHw3vIAuNVa1HSFIUN+bx?869@i+rJ-3s:vN,@v\\\"\\\",2):f(\\\"\\\"}.H7Zv>s+b1b4q+b1s5sk8*s8;CaZtPWcr9ukiDsPWcrvbJt7b4t|8Bs8T\\\"\\\",2):f(\\\"\\\"}bdMAa6*xCvbyr9V@sp1mvL6NvHw5vy<vy5JK*nAyrh.RaR5/vub,\\\"\\\",2):f(\\\"\\\"{y7by+bX\\\"\\\",2):f(\\\"\\\"}UaG/nAU0ib/v9br\\\"\\\",2):f(\\\"\\\"}PaHrRa+EA0M*,beu4.W5njXphv=-/bZacdGNmz6NfDaa8qawCaub|bRa=xm*+tm*Y=ab/bXpn2X>@Bq.C6w.@SWaXI+S,bD=FaO=32L=w*>Xc;c|bhb6CfbqvU|hD,*WaAa,5ozUM|yabo2Fk1wK0BWHZ\\\"\\\",2):f(\\\"\\\"{OJT>=u=OWWa"));
$write("%s",("abhbr*AyL2Sa7=i*f=7b9bsAdyG=Iv+M<av<ubSwQp=>:xQa,bTa.bzbFaP*U1w.B+6bNot\\\"\\\",2):f(\\\"\\\"{fC-ZjUi9gsLpVXITcv8MdbP3+b8r=a7wgM+M<a2b,bubQwY\\\"\\\",2):f(\\\"\\\"}9b6b9bkbi.Xpuyns5w3bZs9b\\\"\\\",2):f(\\\"\\\"}@YQTa,si9ki@+@a6\\\"\\\",2):f(\\\"\\\"{fc:r7b.wFHw-eAfnaM4YGpD+6.*Hyy,FirbGpL59baZT-hbdAqy9-;>Paef+|e8Z<7bHrjVWa.b\\\"\\\",2):f(\\\"\\\"}bp\\\"\\\",2):f(\\\"\\\"}S\\\"\\\",2):f(\\\"\\\"}T4I:9bJ|wtMs\\\"\\\",2):f(\\\"\\\"}bp\\\"\\\",2):f(\\\"\\\"}y>z=\\\"\\\",2):f(\\\"\\\"}b@aGNK59b5bLzE/5OXpU=\\\"\\\",2):f(\\\"\\\"}bq34b7=h\\\"\\\",2):f(\\\"\\\"}i::,xh=3afb\\\"\\\",2):f(\\\"\\\"}QKH6bT@T<z:Vaq:Ooz=@ObR7g6bT@T4|N3,>27/9bbb,b.bfbmbyjtb6bsAQ8Z<7bcbx.c9hbhbc\\\"\\\",2):f(\\\"\\\"{jrQ.K\\\"\\\",2):f(\\\"\\\"}0R@a:yp\\\"\\\",2):f(\\\"\\\"}93a@a>aHra|MEQ8Va*u\\\"\\\",2):f(\\\"\\\"{G;u4bHst<lbC|l9Ua@a;@oL0/+0Aaps8b;r<aTBfBWaW6Defa^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\"));
$write("%s",("\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^32^[2fha\\\"\\\",2):f(\\\"\\\"})3(f\\\"\\\",2):f(\\\"\\\"{#v3mja13(f\\\"\\\",2):f(\\\"\\\"{#,4353(|a3891(f\\\"\\\",2):f(\\\"\\\"{#(ntnirpn\\\"\\\",2):f(\\\"\\\"})4201(f\\\"\\\",2):f(\\\"\\\"{#)~4[~4b^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'dZyzFaEp-b=aoph;ub.bmMf>a1\\\"\\\",2):f(\\\"\\\"}Ewbe8h8oj+b1|cSX8:3Pti*c95btbXaNYu|CCgbc\\\"\\\",2):f(\\\"\\\"}8GogzbkbSwzq|OdM.bwL;y=t?CNa-b,hH,syT+<a5F<C69Cal6i*GCkiH6l07p6Ch+ubFa;Bbx2bTlGvU1.BFG6bxb=aPzKfZaxUjdfb|sL\\\"\\\",2):f(\\\"\\\"{w*vqSFh.xv:2l:|\\\"\\\",2):f(\\\"\\\"}T:y7Zaf-Ba3?oq?a/b=aXa<wMY7j9vZaQwY\\\"\\\",2):f(\\\"\\\"}S9vwSw;6QwY\\\"\\\",2):f(\\\"\\\"}AHDakiZE6?QaPDib.Ed\\\"\\\",2):f(\\\"\\\"{SF,2"));
$write("%s",("Yh6bH3P29b7b+0Wa\\\"\\\",2):f(\\\"\\\"}?4N\\\"\\\",2):f(\\\"\\\"{=DTAa?eUa7N*Ci#chOou+0OoSaq/GoWa5;M2lBHnv\\\"\\\",2):f(\\\"\\\"{iwPakiW,sJXa|mkbLpRmx*cxlyVayYxZ<WPD<p*pi>\\\"\\\",2):f(\\\"\\\"{bu;kbE.|w8wGAr/WaD<6+/OSaR.Q=3biu,zlyJwYaAE0=w==tP.Cz*TOyU31bzrDaGNyboqg\\\"\\\",2):f(\\\"\\\"{mFUua1+\\\"\\\",2):f(\\\"\\\"{RpjbzxtW>.up0b5<q|ml*p\\\"\\\",2):f(\\\"\\\"{b\\\"\\\",2):f(\\\"\\\"{|:ys+5ba1?p=l:x+\\\"\\\",2):f(\\\"\\\"{C79vQ2=TRVol(Waka0bY=XKefwbJ4a:aN/\\\"\\\",2):f(\\\"\\\"{|/CC.,zv\\\"\\\",2):f(\\\"\\\"}z@JzRtiROad3V42.X9.E17dzev:>7|Wa/Jr*-F?>NVMfFbibWrDME44A\\\"\\\",2):f(\\\"\\\"{bgbxbYaCa-Emb9E6.-q@ax*Wv.bf>uq2b|8J-.bH7db3Bp@I\\\"\\\",2):f(\\\"\\\"}iDy?|bwSJLl;hCAfyz|I0sw\\\"\\\",2):f(\\\"\\\"{RweUe7vbYaQaaR\\\"\\\",2):f(\\\"\\\"}b5Gi*u\\\"\\\",2):f(\\\"\\\"}JzW*1wZaos-?kdL1C@f5Y\\\"\\\",2):f(\\\"\\\"{51W;m3ywV-2bn?*r=tGaoYZLK3c,b;@hb;s8ja4oh.3abYafuduDtp\\\"\\\",2):f(\\\"\\\"{Iz5bLz1,iF0"));
$write("%s",("b-<X@k1ar|b1wZa/J69OarTslfAOpUa3t=rdb<+zsldnyaMk;Q-:jjwGMhb;s9y7<jbIAibb=Ta2hnq5GAECa9+1k&6ehd;B1bF|Aw5GswHw\\\"\\\",2):f(\\\"\\\"{8y-izI0Da7<Q:=aPa|mKv2.+rE.7w|bjwfbbp2PjzIgY|Dvog+H/\\\"\\\",2):f(\\\"\\\"{41P57bqiKwm3*Ijb\\\"\\\",2):f(\\\"\\\"}bqF,K8q;23Z+b8bqi5HA2+qWa.C6wScsw3BfJo,l;>aIuUM9Vdz=aEs,Hl4fhTa\\\"\\\",2):f(\\\"\\\"}+2NA-nh<55b1-@5WavbFanh1Q\\\"\\\",2):f(\\\"\\\"}YMDhbY?j2xsabCsMr8jg5776K>aYh32L=I/|Dx2hu@a@hKXU\\\"\\\",2):f(\\\"\\\"{Pad5Aa7bir/bDlL*5bwbv|9bh+QakiMSdFu6hb/CY|opxIaia7b0Gqi;\\\"\\\",2):f(\\\"\\\"}~6e|dtb0b@a:DN|L|,>7?A0=aPqq8z=Rwsqki-KoJybhbzb2\\\"\\\",2):f(\\\"\\\"};vqi=pgsol*HiFG8OB2t.qY0wb6sabCa:CQtbxC>/@K\\\"\\\",2):f(\\\"\\\"{+*\\\"\\\",2):f(\\\"\\\"{bDa:D8\\\"\\\",2):f(\\\"\\\"}0Q.QUa0\\\"\\\",2):f(\\\"\\\"}=t3v2Hv<Va<aFaPDlYBqwbWB*th\\\"\\\",2):f(\\\"\\\"}dvPW8pvb\\\"\\\",2):f(\\\"\\\"{b?VD.t;e/:5fHB2Bai>Kp,bW\\\"\\\",2):f(\\\"\\\"}Dl<w<aw"));
$write("%s",("b<w?aO18>nZ.w=y|bi:>Ki:f-8@ki<<;rU<gN+.nPSaK;VE\\\"\\\",2):f(\\\"\\\"}/H<G-@acb4b\\\"\\\",2):f(\\\"\\\"}Dj18@ow+HSaOBAL:q@acblb.zLr=rj18.RrO18>evbbaMS\\\"\\\",2):f(\\\"\\\"}59bye/(6e|bh*fHB2K;r\\\"\\\",2):f(\\\"\\\"}fHW\\\"\\\",2):f(\\\"\\\"}.dZhaMS\\\"\\\",2):f(\\\"\\\"}fHVEC+zs7bTqcbO,vDOBX44*jb7b4*=v9;vL|\\\"\\\",2):f(\\\"\\\"}rpIh/>IUSFcbQ3IyCu-bKWlx2.yb1Qvb<yeTyb2Wvb\\\"\\\",2):f(\\\"\\\"}@OaUC=avP5xc3e#a/>\\\"\\\",2):f(\\\"\\\"}HhxFvbbL;IE,bw2wb0\\\"\\\",2):f(\\\"\\\"{dpZIf5,bP6a.bSa5gt-s\\\"\\\",2):f(\\\"\\\"{2tAyjpu8Q,\\\"\\\",2):f(\\\"\\\"{bUaSls-bbyS-8gu*blb\\\"\\\",2):f(\\\"\\\"{b<r>aUa0bH\\\"\\\",2):f(\\\"\\\"{WJD/W,sJjb*ti\\\"\\\",2):f(\\\"\\\"{+*GtVo5bfwR?9fuVBBbbpr+*bp+rOprgZICa;vDO0*lxxb>3;vWJZ*hbdv6QCaP*M9f3bclYX@KX0bqyD.EadL2bbL8bu80\\\"\\\",2):f(\\\"\\\"}Hvf\\\"\\\",2):f(\\\"\\\"}9qU9zKab<Y:y5bvbP6U=Ca|Ut?.Ed\\\"\\\",2):f(\\\"\\\"{ZafbmbcyCs1z5bs\\\"\\\",2):f(\\\"\\\"{a>o,o.?axP\\\"\\\",2)"));
$write("%s",(":f(\\\"\\\"{O<xfg*tb\\\"\\\",2):f(\\\"\\\"}qyzxYOJ,z;=+Ta@p2sDa5b:Twb:wwbibQO-vONc>b5bNBDa/AOrOCLrubPtC23VWa<>*qLRF9<+H@dbk<3v=aC>Wvkbccvphj0xoshbDaPDbbk11@8s6zIl14eb@1@gPpC\\\"\\\",2):f(\\\"\\\"{UZlb+r\\\"\\\",2):f(\\\"\\\"}rPaRadb-2A2=9LWQ=pxot*1H>tbPq,pC@q|5pM>An*1\\\"\\\",2):f(\\\"\\\"}r3b&6ebdS\\\"\\\",2):f(\\\"\\\"}Y9Y1/b*blb/b\\\"\\\",2):f(\\\"\\\"{D|bDZlbNY;y9Hbxfbd\\\"\\\",2):f(\\\"\\\"{mXbUhb1|9bjW<Pr6Cp=9.GZak1T6IUtwUWRaGO<=zb,/jbIy<y+|X-rv2.p-SaY\\\"\\\",2):f(\\\"\\\"}IE+-b/xUjbopfcv\\\"\\\",2):f(\\\"\\\"{Hr2pw.5/E4gbW=UZJwzqTastlbDBPWcyh7Ua6q@><aJ03=8pZtdz+.FkVa\\\"\\\",2):f(\\\"\\\"}b*bMD2|0|>adRo\\\"\\\",2):f(\\\"\\\"{nSdrtbd5HruA@JK+@Jhm3hU-W|9M7u6W*bbb:u:|;VL4-bOr/WU+uVtb51oj+bNxI,gZHrNaRppSauaA,5b6bQaDiMr3Yn=xbgB(6ecckbsrbu<+6ty,.N/bMqvb0bNaPD8b,bD6<6hj1q<BgBD+EanrRakraM8s\\\"\\\",2):f(\\\"\\\"{uopCsOa6W+.Fkw*mwwLq;ZbFa?aZrYajbX\\\"\\\",2)"));
$write("%s",(":f(\\\"\\\"}i5Pa8qEwWH6WDFJdYId\\\"\\\",2):f(\\\"\\\"{gs=+CpDvvbC30Rdy|/Kzd2eb0QRPHrb-+bNU0TcopvOBeyI|ouhbubZa\\\"\\\",2):f(\\\"\\\"{Spv/b?S+3clb.bNU0z8\\\"\\\",2):f(\\\"\\\"{ab-Zh.CjW|+b*b1zjbWa077bU41|8>hbt\\\"\\\",2):f(\\\"\\\"{8b+\\\"\\\",2):f(\\\"\\\"{C7hvFuZM=aL*0gdu4pp\\\"\\\",2):f(\\\"\\\"{1z;z077bG04bP\\\"\\\",2):f(\\\"\\\"{?.>;tu=k?.>;0X-qbR~6eY2?Sp?<ahZRa<K<a?+5t>=MFZaFai80+/sLYD6OI6DXautstbb:Xt|>=WId\\\"\\\",2):f(\\\"\\\"}ZxtWcb:s,pO1Ipi:f8R|ir<wDZA0utstgpHZap3v<Dvb8bITouap3vdT?VVZHC\\\"\\\",2):f(\\\"\\\"}Vp|Bv\\\"\\\",2):f(\\\"\\\"{|xbv<<7*bIzw\\\"\\\",2):f(\\\"\\\"}39oh1bvb8b75zt69K+V-bpP8kh3=y:yC7jYui:=xib|ubbQqnp5pM>>-*S>39bv:/>ITmubR=FE|bb2@0/X;OS2b5pRwecu6WMzs1q0sW1J0tbjb8>a\\\"\\\",2):f(\\\"\\\"{GaTVibMH.wXaNa.bTv88kAAX@a:Cjb8bhb:\\\"\\\",2):f(\\\"\\\"{tb7br6l;q;<\\\"\\\",2):f(\\\"\\\"{eyabyb|OxhiuL2MpOBD?/bTaY;Da+rbKA1k+EUFi<wfg|E3b7w;v<ahbhp=+@\\\"\\\""));
$write("%s",(",2):f(\\\"\\\"{Va<k9b|@.E=pUpJY+wGpFAtt?IosWyjb*b>q:u-bKXbbnqBaSlP3x1Fu-ITr|9z/BwCar\\\"\\\",2):f(\\\"\\\"{eUNa/v6Nyrbb5R@a+*NK9btr0o*AexGaRW*b1saRYaHr=awb\\\"\\\",2):f(\\\"\\\"}VQr7<77SK69\\\"\\\",2):f(\\\"\\\"{G|VuP.rhbeXE|vF7SQjh14tC6IgL-Tl:RZa/@6|7bPXOBBL<;GazGWJO03\\\"\\\",2):f(\\\"\\\"{Pa>a5p+MR18t-\\\"\\\",2):f(\\\"\\\"{98D1KVf?IV,bD3?nI@CaPaUajFE|4WLP<pa*J-,bxrHrqqLGXwj9PWOC7C0sMunpibopprH@6WM|hcbusIKCE|N92pd8:vJtcveT.5E6>a9;vFsI.\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"{G<z+M>pswqwM5kiK=vbjbUaybL2+bbb*yt?1bH41FCWU\\\"\\\",2):f(\\\"\\\"{U<jbwb1bzymnu+jbTKIvUTtprS7bYDlbzWSaAGAa3br63b>05bn12*T-rW2bx;2-v9EvwPNa*t5bBu,?vTL4D=h1NwoyDaI+4\\\"\\\",2):f(\\\"\\\"}zt\\\"\\\",2):f(\\\"\\\"{d0h*bYatzLy@g?azrLvki/-/C.bgbWJuA4t*kRTZRP<OTHr95jb+\\\"\\\",2):f(\\\"\\\"{PS\\\"\\\",2):f(\\\"\\\"}bdbr|SxkboOMrTFxb\\\"\\\",2):f(\\\"\\\"}@0bI3s0FHDa:rwbI3Q28T9r+;CtzVfpmQ"));
$write("%s",("HrwbRaXa=ampkp\\\"\\\",2):f(\\\"\\\"{r\\\"\\\",2):f(\\\"\\\"{bzBwK|D\\\"\\\",2):f(\\\"\\\"}b\\\"\\\",2):f(\\\"\\\"{yEEub,*H2m?PaYp5;FU?>PzTFmjeT<Id15,-ufu*D6C5EC.1?=a,b*b>ay-O8XT9+Fadc?pUacbI:PaL:zcUA*b3bBQSat,tbR.GKJvNH>\\\"\\\",2):f(\\\"\\\"}QaYy0b=u0TFaR?6s4\\\"\\\",2):f(\\\"\\\"}O1OaNafbwLnF*qYaD\\\"\\\",2):f(\\\"\\\"}eT@BaHlskbM+\\\"\\\",2):f(\\\"\\\"}RcN335wbx-bDat\\\"\\\",2):f(\\\"\\\"}>ubUZITaL5>AebU<R,,bzbdph+=L|C\\\"\\\",2):f(\\\"\\\"{kl-bQH1ZP2b*+xbR,h1TaZhPaRx?tRaFacNopI\\\"\\\",2):f(\\\"\\\"}|<;z3bQat\\\"\\\",2):f(\\\"\\\"{|5?t<aX;AaD=\\\"\\\",2):f(\\\"\\\"{O|\\\"\\\",2):f(\\\"\\\"}dR39Sa+JGONJA?s\\\"\\\",2):f(\\\"\\\"{ki74b3At/,6s<uIu8F+PFa?hY;\\\"\\\",2):f(\\\"\\\"{O=FprbbA\\\"\\\",2):f(\\\"\\\"}T;\\\"\\\",2):f(\\\"\\\"}?9CXrLS*bX1Nakbz4HPTa*tf6cbIvjPcbGtWaZa>CLSFaHrubYaZzF\\\"\\\",2):f(\\\"\\\"{b2d2h6@apu/@+pab2htbojS+y4RpA25GC|a1jp=IV\\\"\\\",2):f(\\\"\\\"}hvU+Ya+vB|GB?|DBN5dv+b3IO0e8|sT\\\"\\\",2):"));
$write("%s",("f(\\\"\\\"}gp3b25Ay44ExwbZaKR4+Eaxq@Rh*KR8>Q3F2q\\\"\\\",2):f(\\\"\\\"}C|K2lzj|cQpIaQB:@/qMnK:5T,H@-<ebN+AaQu;vCa2|/bQu8\\\"\\\",2):f(\\\"\\\"{Ua,bn\\\"\\\",2):f(\\\"\\\"{J-.phCxH-8\\\"\\\",2):f(\\\"\\\"}HvzOD-.\\\"\\\",2):f(\\\"\\\"{bki?39bx;9bY?9bi*1b*b8*lxTa8b3wD<k2H<Lp1<Rp3OXpJxSl\\\"\\\",2):f(\\\"\\\"{Po6R8B\\\"\\\",2):f(\\\"\\\"{Gz|KbbI|Y/ib>aabxH3bbx=qlbgHebwbtp|babir9r|CNaFabbJzmspx8u@rcbWyEsFB+bLrosZs:j>qr*db,Q3,xbJI@<?wp1x8*b074bB2h+9u\\\"\\\",2):f(\\\"\\\"}Jjb-bL42b>q>aE=L4vbvzbNX;bL8*h\\\"\\\",2):f(\\\"\\\"{TNtb3Op.NHa+L,EautUaYp@?hbQH;x9x>;DaTvi-g?j|iO|sDrq?<aD-rjzrAac*t6gc;M\\\"\\\",2):f(\\\"\\\"}23bHP|bC\\\"\\\",2):f(\\\"\\\"}1bayCa*r7btsh\\\"\\\",2):f(\\\"\\\"}6w>pPtD./@fbdyA-+\\\"\\\",2):f(\\\"\\\"}*M|bU9MthbA\\\"\\\",2):f(\\\"\\\"{kiWNAs*tybxhX;WJC|U,kb*bz3QjPaO36bb\\\"\\\",2):f(\\\"\\\"{@<>v/bWpztR+1b9-lyTazb4bQqEvp2DqLtE>i\\\"\\\",2):f(\\\"\\\"{K6HwtbXtyuQ\\\"\\\",2):f"));
$write("%s",("(\\\"\\\"{4u|Cd5CzD3ibJqm,yb1\\\"\\\",2):f(\\\"\\\"{5>93GoyOSaEcs9:5Ra.b;HvbBwp<zO-b3Apxp@J8L:-<4bNA|b<EL;D=QagB\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"}dBr/,h>-wbAaAabbWJ/Njsq?K+lyH@IE<p8bY/H1rC+6C:pMdbkdS4Kz*M5bDvkb1w-AHr12K;k;6bsI3b|;/bmb,\\\"\\\",2):f(\\\"\\\"}AaVydbE9YrB9ebv?r\\\"\\\",2):f(\\\"\\\"}t?T,wxwy>.B2Q:A1;sYawEP*Q\\\"\\\",2):f(\\\"\\\"{wbgbU9ALGov\\\"\\\",2):f(\\\"\\\"}JFm,qy0uAyi3ohh=X8,smbO9X.m0j=7s5b*bKutMVa>td=wtzb>;jb*Du2lbubf>Z.acAa8q9-tblp7b0bxJvb/bu\\\"\\\",2):f(\\\"\\\"}<aY1m5A1\\\"\\\",2):f(\\\"\\\"{JY9O?v:@n+.Zaeb4bs4wb>D>a5MzbWo:x??C6\\\"\\\",2):f(\\\"\\\"}?FkBlRa<+@aQaw\\\"\\\",2):f(\\\"\\\"}8bcbf\\\"\\\",2):f(\\\"\\\"{YaYrJ,SFzqkb6b/qz.az8p/bd2m*U7Aa+bhqG*78oKUqSnWaZ:/bK\\\"\\\",2):f(\\\"\\\"{yGgbTa\\\"\\\",2):f(\\\"\\\"{<tw0bUamwlbBa/5Qj\\\"\\\",2):f(\\\"\\\"{xW.cbub=a=aRa\\\"\\\",2):f(\\\"\\\"}|n5y|-lFuW\\\"\\\",2):f(\\\"\\\"}|bdb2\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\"));
$write("%s",("\"\\\"}r-vOaQ;=a.b\\\\\\\"\\\"),\\\\n(\\\\\\\"\\\"SaJD9b+\\\"\\\",2):f(\\\"\\\"}Hr6b@ak*\\\"\\\",2):f(\\\"\\\"{bNazqxv=H2\\\"\\\",2):f(\\\"\\\"{yLUa\\\"\\\",2):f(\\\"\\\"{b7h0uG0Iltb>5nhm?\\\"\\\",2):f(\\\"\\\"{x=p1\\\"\\\",2):f(\\\"\\\"{Aay,vbhy6.9fSqhxX*Ga9@Vu.bx89bI/Eq*wy7D.q3\\\"\\\",2):f(\\\"\\\"{bb,@aw*G/Z7uby:+\\\"\\\",2):f(\\\"\\\"}djjb>a@a\\\"\\\",2):f(\\\"\\\"}|5b6*xbP\\\"\\\",2):f(\\\"\\\"}hbKxQaJF:,>->v8@-+I9X-ojmBk=Cae8<aAaWa9C7br*ab/\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{ytb\\\"\\\",2):f(\\\"\\\"{q/49>zrT,Ca9b0bd1=9<aEaNaL2;BlbZhTat-0bxhI,mGmImbZrIuB\\\"\\\",2):f(\\\"\\\"{yH|IibfbFa;H5qgH+bL|irlh1qwbQaFaZatcoJgHopOCCaoj\\\"\\\",2):f(\\\"\\\"}.-zai|HFGprYt6bq<+9Ca5pQa*bTl\\\"\\\",2):f(\\\"\\\"}Ji:YaO,dxLu+\\\"\\\",2):f(\\\"\\\"}eFr\\\"\\\",2):f(\\\"\\\"}mrL2@aiJwbzb|B936/Ua,s>aib*bXa6xVaL:3H<uV,T,tbB.pxo-\\\"\\\",2):f(\\\"\\\"{u148wzz\\\"\\\",2):f(\\\"\\\"{bM27bgBYapxC<8;cyg/4bkbwbhbfwBwzD2..bqi<ajbkb6xnhbrZq"));
$write("%s",("8;7@VaQ@z6DaRahbBaj\\\"\\\",2):f(\\\"\\\"{zb=a1bdb\\\"\\\",2):f(\\\"\\\"{2Pa5b;Bw4b-opzbYatbaHP>XpH39byr9tBapp?a\\\"\\\",2):f(\\\"\\\"{byjw2d-YHBaPcBadb*kh?qCxkoCmG-blwPHFaTB\\\"\\\",2):f(\\\"\\\"}qGzXa<7XyQ,=Hmhr*c3,b-qqsQotblwwbWFwH>aRaEa@aebBafHEpzbmbo1,?L61bBanhhsVan,\\\"\\\",2):f(\\\"\\\"}bL6<aL9NyAn,bV6hbkb=a@tj\\\"\\\",2):f(\\\"\\\"{YoVambubebkbab=tY;.\\\"\\\",2):f(\\\"\\\"{Faoq*2PaprfvWtvbi3W=/bI*<2Sw8rUu/tzbSamh<257vbPaKwRan,F=XaP5?at-7lVag2dr@3?a<:Ra3r=qD-AA>aI+Q=g.I-ibDvcbvstsjbHvKw\\\"\\\",2):f(\\\"\\\"{blx9+WrcbIgI\\\"\\\",2):f(\\\"\\\"}i>gb5bT\\\"\\\",2):f(\\\"\\\"}2bfxdxHrH7/wm,ki=0<a?ac\\\"\\\",2):f(\\\"\\\"}3hX;SaN71\\\"\\\",2):f(\\\"\\\"{8pb=Ya4akGfqoEX;Oa7bCj7bgb?4w,KFVycvTDb\\\"\\\",2):f(\\\"\\\"}6bj,@aDaPawCG,xbebeb/b<EFa,FQE?D,bwbEuvy;7Oj>CsrU<zy8bq4*FWsFiPaVaSnUaT<M?2@Ta\\\"\\\",2):f(\\\"\\\"{uyur6OaAa3Em*CaBy.EQwJ?K5bv@?\\\"\\\",2):f(\\\"\\\"}vAa21c"));
$write("%s",(";T,IE/xOagbZAXamb,b;xvp197b,b1xU<Hr>al8-w>-bbqy?>A\\\"\\\",2):f(\\\"\\\"}h\\\"\\\",2):f(\\\"\\\"{ibaBB9-E\\\"\\\",2):f(\\\"\\\"}bu?-d.E0bc*\\\"\\\",2):f(\\\"\\\"{b7?=aOAtnasYa+4Dae-CsXaE9*veb/zEvVaAaWz8bh\\\"\\\",2):f(\\\"\\\"{dzArGab6,bKuY\\\"\\\",2):f(\\\"\\\"}W\\\"\\\",2):f(\\\"\\\"}?a<aub1ba*.6fx\\\"\\\",2):f(\\\"\\\"{qGz9.o4nwo4vkmEB*mCCCwbNxXa\\\"\\\",2):f(\\\"\\\"{bol9:5<\\\"\\\",2):f(\\\"\\\"{x|;@ss:mrXau|C,>5WaB\\\"\\\",2):f(\\\"\\\"{m;BavbhbW;5|U2v1QuNaA9Na\\\"\\\",2):f(\\\"\\\"{3>9Y944Yh4;z;bBfb+z.6-bOAFamh,\\\"\\\",2):f(\\\"\\\"}h,tbyuPjA1Bf,Dw\\\"\\\",2):f(\\\"\\\"}r.>q1bVaXt3bUaRambVaZaNolbHrP3fu\\\"\\\",2):f(\\\"\\\"{2zqn1Dth,Yay\\\"\\\",2):f(\\\"\\\"{olh1k2X;mbGxUac*x=aD3s;,A4?Ckpd|Ya-biu8yHrcb69,bW2>aT+vb8;Tx@aV-13\\\"\\\",2):f(\\\"\\\"}q0b6bo4f2l0+bhb\\\"\\\",2):f(\\\"\\\"{|L:kbPa+b6bTakbxbZa>1m*-b,B6bHrCzc*+x\\\"\\\",2):f(\\\"\\\"{|Lu2bz:Qcdx5b9?+bE+3/j|R<D:E*jA*khACa|bC3ab8bMpOaY34bKf"));
$write("%s",("ryMuXaq-krfhw.L9?aw,=wF3==abxbK>Pa.bY/FuXsgY2btbZ.gbX7jbhw/bWamj:8yb@a;s:iD+ymIzDis+0b<a\\\"\\\",2):f(\\\"\\\"}qC3Iz4bG+fh1bH\\\"\\\",2):f(\\\"\\\"{Y/08lrxbY.EpU*n,@6P6bko1m;Qul2j2SaNaeb\\\"\\\",2):f(\\\"\\\"{bs.v.WaEas8.q2r@a|bgbQwr.ybOar.P3FaNp8?Ig?abbHr:sR5mbOa9rkb|bs\\\"\\\",2):f(\\\"\\\"{V8R?<*zbL28>Aavt6vf1Xq4bdbWa+.QzEa|b,\\\"\\\",2):f(\\\"\\\"{vs6b-bjd:iybxr\\\"\\\",2):f(\\\"\\\"}bX.e9VyL@;@Eaw\\\"\\\",2):f(\\\"\\\"}U7bb;@YaX.7/A4lb.bj|582ye?\\\"\\\",2):f(\\\"\\\"{kc?9bPa>;55J@H@D-v8kh4b\\\"\\\",2):f(\\\"\\\"}bQaAiHr9-F\\\"\\\",2):f(\\\"\\\"{3bM-WaT40/?ae84@kbgb9;5bkbx2>aGaQ*U*B<X8\\\"\\\",2):f(\\\"\\\"{z7bybki+@lbZ*3bl1az:y7bmbkbFalv\\\"\\\",2):f(\\\"\\\"}bHri\\\"\\\",2):f(\\\"\\\"{M+hb4bl18bHx4bt6x;\\\"\\\",2):f(\\\"\\\"{vHn\\\"\\\",2):f(\\\"\\\"}r1q5.dbc5l@Pwh8h7\\\"\\\",2):f(\\\"\\\"{>=,c2Euey;<5|<a1bFqi94bUrs\\\"\\\",2):f(\\\"\\\"{L|Xpquo1bbirNp:9n?tb0*Z.ubx>mz1rH9*;kbr>U7kbA"));
$write("%s",("ajbCu1rxb2.DavbAaib8bM>5b,b4;d\\\"\\\",2):f(\\\"\\\"{/5T\\\"\\\",2):f(\\\"\\\"}BaQa|bw.IvXa6b<aibG|m;p\\\"\\\",2):f(\\\"\\\"{z<x</b<9VaBaNamhabSa|+2;4t\\\"\\\",2):f(\\\"\\\"{k@*Q<*kO<H1M<Mpc+|blhjbU*r\\\"\\\",2):f(\\\"\\\"}@aPaYa=1>aYa4,13jb1b2b5b\\\"\\\",2):f(\\\"\\\"}wgzzbx8Ta51Fa\\\"\\\",2):f(\\\"\\\"}bS|AambDaNaVq=adb-qzbC,ZtAr2tb=N,mnkb8bL6,q-1+bTrg.91T\\\"\\\",2):f(\\\"\\\"{;|j\\\"\\\",2):f(\\\"\\\"{usnp1rRu1rX9CagbD+WaV-B+0+|bYgDai\\\"\\\",2):f(\\\"\\\"{Zq-bx8ubXqY=Oar\\\"\\\",2):f(\\\"\\\"}9bU=ZaD+1bEp+bDawb5vm*3bB|33vbp.y87b\\\"\\\",2):f(\\\"\\\"}b,b3bHrm22b6xibr*Ya3b6bdbRaNaI/Vau4@tu=jbzs=6VaXsi3@ahv/vWaC<AaOa.b/;=aWa694b>aw,+qIs/b*\\\"\\\",2):f(\\\"\\\"}=aEaZ+QaEaM2Oam3HrjrVaZhtbVa?aQ6;zL.C.8b3bTvm|G1\\\"\\\",2):f(\\\"\\\"{kC*j|A:=r1.o0X8Sau4mbUaAaSaVaD-1qWv2*Hr3bwbCagcryXa=10b3p>xt:\\\"\\\",2):f(\\\"\\\"{bE+olRwjbq*2bywU0=aq8ibBah1d0,bG/lb:rybdbhxDv5v<;YrBa0bf*"));
$write("%s",("C\\\"\\\",2):f(\\\"\\\"{xp.q\\\"\\\",2):f(\\\"\\\"}s=|7;:j.xztQa4bub5sNhIzAaj63bU013\\\"\\\",2):f(\\\"\\\"{zzqlb+b3b1xX8yr5*Yr8b0bj\\\"\\\",2):f(\\\"\\\"{O3YzWzgbqxTaebf/7bRaTaIvUaEakxz+AyUaTa\\\"\\\",2):f(\\\"\\\"}b5,Ey1babovCa0hQaZzkb<*J-Uatb-ur|4bRa\\\"\\\",2):f(\\\"\\\"}vXa.bXawwDl?rR1ibdb4bisfk<r+\\\"\\\",2):f(\\\"\\\"}Xalp2*-b-h,b\\\"\\\",2):f(\\\"\\\"{b7ljb/b4bNaXa3b@a\\\"\\\",2):f(\\\"\\\"}0g\\\"\\\",2):f(\\\"\\\"{Ra?vPahq,6?/F168|6Tr:sRaV-ybXpcrlb3r94Lyi895bb\\\"\\\",2):f(\\\"\\\"}u\\\"\\\",2):f(\\\"\\\"}v3b|uzuWuUt7\\\"\\\",2):f(\\\"\\\"{jbXtb9,\\\"\\\",2):f(\\\"\\\"}gbvb,\\\"\\\",2):f(\\\"\\\"}QaecSqbbZy:vVal4b\\\"\\\",2):f(\\\"\\\"{xjJt4bbb/bUaQ,z,H9B\\\"\\\",2):f(\\\"\\\"}azebNas8Z.kb\\\"\\\",2):f(\\\"\\\"}b\\\"\\\",2):f(\\\"\\\"}bPamb=ahb@aAaohBaxbVtzb*\\\"\\\",2):f(\\\"\\\"}1rDaibCvbb\\\"\\\",2):f(\\\"\\\"}babdvr3hwc,Ask/XaxbIv8s9g\\\"\\\",2):f(\\\"\\\"{tPzOa*bYtfbEpUa>adx9bCt*bFar9ap4b,bUqZaRxBaHr\\\"\\\",2):f(\\\"\\\"{"));
$write("%s",("y?a6byblu6ps3/b<a9bFa0bDa\\\"\\\",2):f(\\\"\\\"}q\\\"\\\",2):f(\\\"\\\"{v\\\"\\\",2):f(\\\"\\\"}bfbZzzjTaoz@-h1lb\\\"\\\",2):f(\\\"\\\"}b\\\"\\\",2):f(\\\"\\\"{*xbI|nhUae8hb-bJ,r\\\"\\\",2):f(\\\"\\\"}d,Da7b=a\\\"\\\",2):f(\\\"\\\"}q8bq8BanjU7u6SaFkDaz8uyw8\\\"\\\",2):f(\\\"\\\"{byphqQv48h4dt*6Fc<a-u-bfvkx5b1bOaDqevK\\\"\\\",2):f(\\\"\\\"{?a9bdy>aRmibFadb\\\"\\\",2):f(\\\"\\\"{bv7\\\"\\\",2):f(\\\"\\\"}bA7kbtbh*fb0bFuwblbR,2gubOaKzopybNacr.b*b\\\"\\\",2):f(\\\"\\\"}bgbM-bbbbfc+r55\\\"\\\",2):f(\\\"\\\"{b>aq.ablzolUaC\\\"\\\",2):f(\\\"\\\"{-.4+2\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{bwb8ro737qqN5+blb-.53B5hbo\\\"\\\",2):f(\\\"\\\"{o7Vaubfctblz:s1sk7q6brV,|-azopDvubRaQ\\\"\\\",2):f(\\\"\\\"{:5/z50ebjbxbg.6blb1shbevx2cj>aJw7,yb<aBawb1q\\\"\\\",2):f(\\\"\\\"{jA0=-C,cbJoAab5UambHrP1-zi\\\"\\\",2):f(\\\"\\\"{,bC6DyT,YadbazFaabmbi*F2=aqy=y.bYa.bo2;\\\"\\\",2):f(\\\"\\\"}@a:54xVoa.Yaxb6b7*LzZa9mH13y>/j-i4lb8bz.Hr\\\"\\\",2):"));
$write("%s",("f(\\\"\\\"{v9zybUa4e7bSam\\\"\\\",2):f(\\\"\\\"{.b+tJuzbCaTafbjdXqgbxu0hkimm7zHrGav/mbxb12=yWa+bQaxb4sNaYa,b2byb>,o*r|kuw\\\"\\\",2):f(\\\"\\\"{bbZtVxi.?aB\\\"\\\",2):f(\\\"\\\"{ybPabbBaab7bIxWrB+3b7\\\"\\\",2):f(\\\"\\\"{ec?nmb:xcbAa\\\"\\\",2):f(\\\"\\\"{.=aSaQ.2.QaL46b2bHre-ms5zypOa5s32cy5b4b*b8q2bJ\\\"\\\",2):f(\\\"\\\"}Wap\\\"\\\",2):f(\\\"\\\"{kbQaCsDaebZa2s=alb7bZ0K3eyEafb\\\"\\\",2):f(\\\"\\\"}vs1cb+4CaQa8b-vcb5sub5qozHrJ\\\"\\\",2):f(\\\"\\\"{W1LrTaPahbCaRxl,wb3vdbEs1bK\\\"\\\",2):f(\\\"\\\"}CsjbPa*bSawyvbeb<aFgibl1ZxW\\\"\\\",2):f(\\\"\\\"}KwubxpYvFaEaSawby-W36bbcQaQaTaCaFgVvf4/yI1C1EsOshbabdbo-kbxvm\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"}bRa;1Xvu0*bmbCavyvpv.4.YqabFacb3b3b5b\\\"\\\",2):f(\\\"\\\"{bEaZrHrzb/bBafb9b*bkbLr.bkx*bgkHr+bdbKqS0xbvyUuUap\\\"\\\",2):f(\\\"\\\"{G02b7bSoqyR+vbNa8qe/dpEa9bY.8bi*vbEaibyrTayb\\\"\\\",2):f(\\\"\\\"{|*b9bBaWa*b5\\\"\\\",2):f(\\\"\\\"}f*:zUzr"));
$write("%s",("g6utbBaL\\\"\\\",2):f(\\\"\\\"{R,lbib/,IyVaQakbJzbx>ah.,bp1C|RpcbxbQaQuD\\\"\\\",2):f(\\\"\\\"}12>aRuki.2,2*2-v\\\"\\\",2):f(\\\"\\\"{2Cj*bco\\\"\\\",2):f(\\\"\\\"}bSuT,JvPa6b8bFa6b/\\\"\\\",2):f(\\\"\\\"{*bnjwbvb?aJ\\\"\\\",2):f(\\\"\\\"}5bEx4bP0N0ibOaFakb3bXaC\\\"\\\",2):f(\\\"\\\"{ib*|4b@as1fb3bhbYaPa2bAaPaD\\\"\\\",2):f(\\\"\\\"}mbPai\\\"\\\",2):f(\\\"\\\"{BaWvSaBa=xy|fbWahqUvm-;/Tv=/yik-,wab\\\"\\\",2):f(\\\"\\\"{bJz+bWa0o0b51Ya6.4.g.lb*|GuXafh./J0+\\\"\\\",2):f(\\\"\\\"}FaJvI+tbFr8\\\"\\\",2):f(\\\"\\\"{xu6ze|c|3|1|+rKz?aTaMotbab4bcoPafbBahpmbmbtb@g>aU0xxBabb-bT\\\"\\\",2):f(\\\"\\\"}/\\\"\\\",2):f(\\\"\\\"{ksYa8bCaqv6*dbmb*b-,vbdbdbebt,cb+d>0Wa2b>aebfb,\\\"\\\",2):f(\\\"\\\"}Hr|bco+0\\\"\\\",2):f(\\\"\\\"}b.09b.09rRa-0.0+*+0?akb+0UaUqWa-bjbB-Uq./CvHxnyQ.ab+\\\"\\\",2):f(\\\"\\\"{o.Ua6nUq?avpUaOaS/f/f0Q/O/P/I/lbG/WaAu*|kbbbYmK.S/L/hbP.K/Sai/*bRai/<af//bUqQaOa0/kiJr7/hq</it:/Rvj|F*hq"));
$write("%s",("dd+\\\"\\\",2):f(\\\"\\\"{Ra4bzb0bRaDzlbgbWa1bSrh\\\"\\\",2):f(\\\"\\\"}Vab/Eagbq.o.t/u/kis/q/HrDaVaRa<aWaUq,b+*Qa=a\\\"\\\",2):f(\\\"\\\"{bRaSa=a+b?aSa?ambXaUa3bDalbVa.b@a.bRa=a<x2*Balbj\\\"\\\",2):f(\\\"\\\"{1hppEaAaHv+b@aSa>ai.-x8bmb=w4bwbTqmbYamb\\\"\\\",2):f(\\\"\\\"{bWaXaXuEax.mb@appOay.CaSa.bTqWaVaSaWakb.b*tabXaZa.bZaabryUsjx\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"}Mo1bcbvbOa6xBy8qvzgbZaCy-b4rOa>aSa.px-6b5u*b6bNa@a9w*bSoBaAadb/vOaUqOoVacbIytbRam*Eq8bWaTiAahvX\\\"\\\",2):f(\\\"\\\"}JzgbPaDa3w2bVaUav-gbouy\\\"\\\",2):f(\\\"\\\"},bK+3rzbRargK+\\\"\\\",2):f(\\\"\\\"}q5b/b>,Wajb0byiD*5yh-etqo?*0hCaVaFaQ\\\"\\\",2):f(\\\"\\\"{ubJuX\\\"\\\",2):f(\\\"\\\"}SaHr8bibtbHr5gFavbt*tbQa6s0bly<aebUaibQadb:,,bQozb;*5\\\"\\\",2):f(\\\"\\\"{ebYa|xQa3bebRafbExcb?xlbPa|bxsZadyzq@aI|XaOaol<aUa/b4w8b@ggp=w\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}Ktw*4bYaDaubWaSjKzfbbbAy,bPaNa2b1"));
$write("%s",("bkdSa-qjwbbQafbPaCambzb=tzrlbkbouZakr1blb\\\"\\\",2):f(\\\"\\\"{|<+kb7bzb@a3w*b*bdxzb<a3wv\\\"\\\",2):f(\\\"\\\"{-bi*1lkiq+lb;s3bMufb8\\\"\\\",2):f(\\\"\\\"}qyVtN*ZaSacbI*-q0b/bubtbQz\\\"\\\",2):f(\\\"\\\"}qTabb=z0bPziuZa1b@tEat\\\"\\\",2):f(\\\"\\\"}Ta0bKxTs=qzx\\\"\\\",2):f(\\\"\\\"}vK\\\"\\\",2):f(\\\"\\\"{Qu>aZaYa+bM*Tawbp*kiImkb-hWvhb>adbEaub9mTviovkA*0y\\\"\\\",2):f(\\\"\\\"{ih|i|l|-qRw.dMt6bBp|bDrVaXa0bOaXaPa\\\"\\\",2):f(\\\"\\\"}b2rbpgbUalbCrybCa\\\"\\\",2):f(\\\"\\\"}brjHgvbVa.\\\"\\\",2):f(\\\"\\\"{DafbkbTa?xZa5b\\\"\\\",2):f(\\\"\\\"}sBaTa2bOa0bfbZa8b|bYakb2\\\"\\\",2):f(\\\"\\\"{SaXpmbBacb*b=aYaRaCzt\\\"\\\",2):f(\\\"\\\"{xbEa0bMpqvOrcbOawbqszbC|2bYaNa\\\"\\\",2):f(\\\"\\\"{bZbzqPaXayr|bdpvb<ad\\\"\\\",2):f(\\\"\\\"}vs-bZa6bcb+r*bAahhCjjbTaUawbEadbkp-bDq.bPa3bZa>leb|b2bcbu|psNa+uCaY2f\\\"\\\",2):f(\\\"\\\"}=anw8b7xFa7bhbWacb6bYaub+\\\"\\\",2):f(\\\"\\\"{9bcbabQa5bQuFaMscb.b+q/bEaJwXa"));
$write("%s",("7b2bQu*b+bgbC\\\"\\\",2):f(\\\"\\\"{mb\\\"\\\",2):f(\\\"\\\"{q*bEaYaSwcw|ywb*bdbNaB\\\"\\\",2):f(\\\"\\\"{/babBaSz\\\"\\\",2):f(\\\"\\\"}bMxbc>awb,by|NaegUaNuRabbNaRttbPawbEtYvhq|kg|Ib6y.yyi,y\\\"\\\",2):f(\\\"\\\"{bOadbvb5xab,bhbApXqjbZa,b5xYqRa=kWy6u\\\"\\\",2):f(\\\"\\\"}rwbNaOaPaxbYyVaUiXvtbcbCaybkb|q6bhb3b0bOhdbkb0b?a,b>a-b+bZa|bWaubab1bQaKt4bhbYpxbAa.bDagrAaabWahj,bFaRpfb/z-z8bAaFa/bAa1wDaWalbCa3bmbEambqtZasz2bSwVakb*z|zzz8bwbUabbfbXa-v=aOaTaAa1q|bhyAyHrlbWa?xkb.hcbib5bYp,x>afbibwbXaRakbVaZribVaYaVabb6bQu3bSafbabTahvXx/bJpgb0bHr,bUaXaDaCjCv/b=weu\\\"\\\",2):f(\\\"\\\"{bXa@a*bOamb6b>aRohyolHr7p,b;vdb0b3vAaXa,bibEaAfib3bCaWthvpvmb-b-b\\\"\\\",2):f(\\\"\\\"}bDaRxyi4ykt1yjqht-yftTvlqvkSvFrrrhu0bZawbebCaeb8b7bnyPs1bPaFu>aNalbwbKuSudvibfkcb8b/bXaeb-b3bZqfvdv\\\"\\\",2):f(\\\"\\\"}bMu3v4tHrSpJtFr?aab9ivbbbmb4b:i5bYafblb?a1b@sS"));
$write("%s",("a+rwbPaFamb5b=aCadb=a3bOaab|b/bPa0b8b+bRa+bupSj\\\"\\\",2):f(\\\"\\\"}bSauf7b\\\"\\\",2):f(\\\"\\\"{bCa.b,bybmbAa\\\"\\\",2):f(\\\"\\\"{bZt,p\\\"\\\",2):f(\\\"\\\"{lub0b+bPtwb6rlbjbOaLslbOhdrQr0b,tWp@i<w0bmbebFamn8rpukwibjbEatbwq?r\\\"\\\",2):f(\\\"\\\"{b4ryb.bmbabcb7bXaQaqs,s6b\\\"\\\",2):f(\\\"\\\"}wYaebEa?aHryw/bdb7bZa0bXa\\\"\\\",2):f(\\\"\\\"}b+bYabbGvFk\\\"\\\",2):f(\\\"\\\"{b+bibHrmbwbub9b|bNaCa7b7bMq?rmb7bfbIoBagbvf4p6pbb7b.bebib9m4altPvlohqctbbib2bjbdbcbSa6b\\\"\\\",2):f(\\\"\\\"{b0b\\\"\\\",2):f(\\\"\\\"{bubdbztcs1pdb,bSadb5b3bEaVapugbmbGa<sUuWaSaTa6bZadb@atb\\\"\\\",2):f(\\\"\\\"}b8bOazqzbOa<atr,b4uMu0beb\\\"\\\",2):f(\\\"\\\"}bEaQuubAa>a\\\"\\\",2):f(\\\"\\\"{bCjYaYqSaubgb1bbb4uvbcb-qwueb5b>aQatbgb*s4u@a-bhbgb\\\"\\\",2):f(\\\"\\\"{bAaDuub7btbdb*bebHrSaSa|bkbHr9bvb,bRa7bNaValbbb5s-bYaolZtOaQo?a3bTacbmb3bcbfbUa5pebTa<kRa5bNazbfbvb1bubNa\\\"\\\",2):f(\\\"\\\"}bVa"));
$write("%s",("tbfb8b5bjbCa+b\\\"\\\",2):f(\\\"\\\"}bjbubibib4bHryblbTagbZbSrVajb,bHr,s*s4b+bTaZazbyt>rkbWa@aUaLr,b.p@g|bFrTa\\\"\\\",2):f(\\\"\\\"{b-b*bfbzbSrvbTa@fFrYalb9b1plpNa@rbsVa5bRaBa8bgb4b=a@aLoyijtdqgtoo,mkqgqhq<maqcbQaUaGoabzbWazq3bibmj\\\"\\\",2):f(\\\"\\\"}bNadbOa/boqnpSaEaHrfhubHr\\\"\\\",2):f(\\\"\\\"}b6b7bdbwb2bBakiGrOaxbBambSa0bPa?aUa1bFa.bibmsgbQa1bfbOa8bUaQaSc,bjp.bTaQa>pfsSa9b2bFaebOa1b5bcb<a7bkb5bAr?r=rSaabubjbcb9bzbjbRazb2b:rebjdQa9bHr@aGavr-b\\\"\\\",2):f(\\\"\\\"{b8b4b5bOaubQa\\\"\\\",2):f(\\\"\\\"{b.bUaab.b1bkbcbprnr?n?aPaibTa>qjbjbLhPqFa-bEa8bPa,bWaxbkiqbdb1b-bab5bDaYaQjDaUaPa7bDanh1bEaEaFaxbcbYaabvb@aublbRa@awbLhWaBakb+dXayq*bBauqtccbTa,bvbubCatb2bdbTatblh3bAa0bdbCa>a,b@aNa|bAanpmb0bcbOh>akbNa4bXabbhbNaBaDa0bLhhbwbdbDakbvbhqko\\\"\\\",2):f(\\\"\\\"{ibq:meqmoyicq/mpozkno3hZakbebJp5b\\\"\\\",2):f(\\\"\\\"}b2"));
$write("%s",("bCa5bmb\\\"\\\",2):f(\\\"\\\"}bcbwbabDaFa\\\"\\\",2):f(\\\"\\\"{b7pebegkbdb+bOabbablbmb>agbBa2bTa-b6bib,bdb\\\"\\\",2):f(\\\"\\\"}b.b?aDaPoCaabwb6b/bypzpxpvpgb7b/bYavbDaopRaRa>aFa|bebzbdb8b<keblbzb,bNa7bvbCaEahb<aCabb*b8hQaub*bWaQagbSa,bEa7b6bAaEaUm>ofn*owouoXf*o*n?aSg4o;a2n\\\"\\\",2):f(\\\"\\\"}nuo\\\"\\\",2):f(\\\"\\\"}oQm.o-b*o1nCa/nWnwbic8aZnEnFmxoEaQmFntn-a8npnnn9m\\\"\\\",2):f(\\\"\\\"{ijo;mho9a9m*k*k-m9m/b\\\"\\\",2):f(\\\"\\\"{f-a;hub@h|eQnIn<nMnDm9aEaOa>mvnGm/nVmzn2i:a>n=aAa/n;nCafnwn-n@a<a-b2n6nWm2nYmEm.n1nAa:aCa8a+n>aXmPmenZmKmhnAa0lWm|eqnzbHmbnImSmBaEmOmMm*bvbtb/b-aJdHd>manRmWmUmSe|eNmTm?aAa-aDm8aJmHmFa@aEm\\\"\\\",2):f(\\\"\\\"{bCmHaAm9a|eBmxb8a+e-a1beg>mum8arb8aXf9m9mMi+k0m6l@l,k7e,j*jokyi.mvk+myk\\\"\\\",2):f(\\\"\\\"{i\\\"\\\",2):f(\\\"\\\"}knm*j6b-a+czbxbubHaqb6aqbEiFiDi5aqbebYi,bAfzb.bKfnbxb\\\"\\\",2):f(\\\"\\\"}ikiZgXgag"));
$write("%s",("IkAl2j.kel?a=aLi;dLf7lRi5luh3ltcBa3aPhIgDiwbPf?aRkYkNkBa?aKi6e;hrbTk?a7iQkvhOkDa?a>aKi2b3bGiUfTj8f2i-b:kCa3aKa\\\"\\\",2):f(\\\"\\\"{b;a3gwbccIa3b1bbk,b|b0auh\\\"\\\",2):f(\\\"\\\"}h6hlk1jjkCaKi.bti0kkkMi.jyb3bKk7hDh/k*h-kBaLiMf1i\\\"\\\",2):f(\\\"\\\"{g\\\"\\\",2):f(\\\"\\\"{gsbubwbki-a;k9k:a;b6k1b0b-b3aAa3a7b-aki.a:b:b,b?a3j5i5h0jik4axi\\\"\\\",2):f(\\\"\\\"{k\\\"\\\",2):f(\\\"\\\"{kwk3aLiyiuk-fzi-j5e+jmdrjRf7hvhQiOi/j3a;hwb+b-aPcPj/b8b1bPcxb;aUf-b:fZapg|b.b5b-aHj>i3bWfvb|bIgGipgfg3bgf;a<b:b3b-a8bIg,bxb2b2btb;a7hWhPimiNi@aKiIhujxbsjqjabVaTaRaOaHa6eEfOhFfjb-agbebbbcbZaVa-abbVaEf-aZabbebSaHa@g-a3hhbQabbZa7h*h6iPa4i3a>a3a5anb-aEi/b3b4b.bHa8byb2b2gtbWfxb5b+bYg7h5hliYhWh;d+cKfHa-i-iFaGaji|fld4a.gwi/auh4a-afgdgMaFa=aWh-bYhDhChGa+bJdRh9a\\\\\\\"\\\"),\\\\n(\\\\\\\"\\\"/b5a|fCc8g-bPaBaobDhHfMa9aMaIa5axb3b.b4b0bxbzb-btbeg7"));
$write("%s",("hkg5hGaMbHg2bzb;azbLfccJa7b?a?auh*hCdYaOaVafbVaibNa=avhvh?a;aSgVaNaUa.guhkgvbpbEa*c7b@aFaDaDa>anbJdubSczbPfIcQgyfwfuf2bsfNd3bHa?e-a-fZf:aIa+c9f:avbldub4bcb-b3ggc0gHaebdbJaGagfef8a1bxbwbtbxbUaac|b3bdgfb/akgzgtbxcRf?a1akg-a6a5bhg>azd:a,cNahgwb.b;b>aagob,c:a-a.b\\\"\\\",2):f(\\\"\\\"{bvbxb5a1aob,fCe2b-a:b1dtbHa6a/c2b/a,fPcFf/b:b6aKa6e1b4eIa8btb1b1bNaGatb5a+ctb,b-a\\\"\\\",2):f(\\\"\\\"{fyb3dMd-aDdBd@dmf/aob5a.d,d*d-b4b7eSc;axb+b.bbcZb0cbfJasdHa/aed+e0cGb/d,btb-b4aWbudpcgdLc=chchd6areOapc0cNb/a;bje/eGaHb5dedOb.a8aNd8aLdLa=a>aIaOaJapb6a+e5azb+cdcfbhc;aOaFdYd6aHaCa@aIaQd8aHa=a.cIbCbMd\\\"\\\",2):f(\\\"\\\"{cycvcocRapcXbocTa;b;bpbgbYdJaGbRanbQaJagbnbcb>dqc5dpbebnbOa8a0c4aJaTa5a+btb5bxbJaQa,c*cRa5a1bzc6aedMa0c3bldjd;aeded8ard5a6a5aedxb/btbvb2bxb,c1b4b3bxb1b0cocPa8aNapcMagdUc3b|b+b/b2b4a"));
$write("%s",("rcFbnc4a=a?axbtc4aSbJcPbKckcic+bZb3b-bzcXbqcFb5aMa/ancvc+b+b|byb4a9cVbNa5aRb7cFbnbFbMapb2c.aMaFb.=ba4a5aJaOa-a-b|b-aeb5aicybHa<b/akc>a>aXb6aOb/a8a6a/apb4a1b.b3bvb4b1b3b2b-b.bvb4anb/aJaPa5a8a4a6apbEb5a5aBb,b9a4apbpbnb8anb4aGa=a:bJacb!\\\"\\\",2):f(\\\"\\\"})46(f\\\"\\\",2):f(\\\"\\\"{#~[2xha=s,y=z,13&X3^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'yay,]99999[gnirtS wen=][c n3aea\\\"\\\",2):f(\\\"\\\"{)v]y3b&a(niam diov citats cilbup\\\"\\\",2):f(\\\"\\\"{RQ ssalcz4rfa cdlnl3c/a;maertStnirP/oi/avajL tuo/metsyS/gnal/avajm4bdateg@3doa2 kcats timil.v3dga]; V);Q4aC3ecaL[b5aX4hha dohtem?3e;4nga repus&3ecaRQ@3cgassalc.<"));
$write("%s",("5joa(=:s;0=:c=:i;)|4ajaerudecorp/3fqa(tnirp.biL.oken\\\"\\\",2):f(\\\"\\\"{.3bianoitcnufR6\\\"\\\",2):f(\\\"\\\"{sa(rtStup=niam^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^32^[2fha\\\"\\\",2):f(\\\"\\\"})3(f\\\"\\\",2):f(\\\"\\\"{#v3mja13(f\\\"\\\",2):f(\\\"\\\"{#,4353(ga36(f\\\"\\\",2):f(\\\"\\\"{#j4[j4boa(etirw.z;)tuo.N8aba(67b~auptuOPIZG.piz.litu.avaj wen=zG4Zka91361(f\\\"\\\",2):f(\\\"\\\"{#tm4[m4c5aR0Z0Z/512152353/2/2166263=4/3141726??:1518191:1/@4[@4cda*6 Q5[p4dea1312^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\"));
$write("%s",("\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'5[w8[$5ofa41310r4[r4c7=[B>[j4[^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'6pma(amirpmi oicy4[(5[j4hma++]371[]591[?6[?6cpani;RQ omtirogla\\\"\\\",2):f(\\\"\\\"{4[\\\"\\\",2):f(\\\"\\\"{4cua;t:\\\"\\\",2):f(\\\"\\\"}%%%%\\\"\\\",2):f(\\\"\\\"}fi\\\"\\\",2):f(\\\"\\\"}*-84\\\"\\\",2):f(\\\"\\\"})48z3b(a]i[\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"}+17\\\"\\\",2):f(\\\"\\\"{<84.;i:-i602\\\"\\\",2):f(\\\"\\\"{;i:911\\\"\\\",2):f(\\\"\\\"{;j:632N4Zsa7218(f\\\"\\\",2):f(\\\"\\\"{#(tnirP.tmfIIcfacnuf;&4[&4bdatmfn4[n4cgaropmi;ILagaga"));
$write("%s",("kcap~4Zea1304T6dbapD6[r4cba-l4[l4bjatnirp tesY>[ca89&AafantnirK7[ia959(f\\\"\\\",2):f(\\\"\\\"{#fp4[ga^64^\\\"\\\",2):f(\\\"\\\"})74[8awa,s(llAetirW;)(resUtxeT:Paca=:R6[ba1Q6ak8ap4[p4adaS Cn4[vEaca&(z5[z5aba 06[06[06piaRQ margo^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'5[t4cjaS D : ; R-5[%L[j4[j4o%6[k4aqa. EPYT B C : ; Az4[56[j4[j4nka)*,*(ETIRW/6[J7chaA B : ;s4[s4aba [2cr4[*5dia: ^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):"));
$write("%s",("f(\\\"\\\"' ohce4B[ka3(f\\\"\\\",2):f(\\\"\\\"{#(stup;Rcdatniy4/ca0153.ea%%%%m4[m4[53ipaparwyyon noitpoz4023[230ca(nVO.ba5FQa\\\"\\\",2):f(\\\"\\\"{aetirwf:oin\\\"\\\",2):f(\\\"\\\"})8(f\\\"\\\",2):f(\\\"\\\"{#>-)_(niamp3c\\\"\\\",2):f(\\\"\\\"{P)ka(f\\\"\\\",2):f(\\\"\\\"{# cnirp/L)l;eja.OI[p]^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'[(3rba@~Wa7;alaM dohtem06x*3c|5aV;cpadiov;oidts.dts &Ya;6n+4d\\\"\\\",2):f(\\\"\\"));
$write("%s",("\"{3kkaenil-etirw~5dva(,^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'s%^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'(gol.elosnoc;)^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'73g\\\"\\\",2):f(\\\"\\\"}a^129^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\"));
$write("%s",("\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"' nioj.)1+n(yarrA>-)n(=fI3cwa^31^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",2):f(\\\"\\\"}54,1\\\"\\\",2):f(\\\"\\\"{.^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"# qes-er()|3cH3bba^31^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"p3lg3fw3hla1% ecalper.j4dea^128^+Ac/arts(# pam(]YALPSID^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\"));
$write("%s",("\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\".NOISIVID ERUDECORPA3cma.RQ .DI-MARGv3g53d|bNOITACIFITNEDI^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"[tac-yzal(s[qesod(^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"))System.Console.Write($^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"Put caffeine \\\"\\\",2):f(\\\"\\\"{(int)c\\\"\\\",2):f(\\\"\\\"} into the mixing bowl.^64^n^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");M3pva^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"Liquify contents of"));
$write("%s",("E3oeaPour^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'3w^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'4e\\\"\\\",2):f(\\\"\\\"{abaking dish.^64^n^64^nServes 164cma\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}^31^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");\\\"\\\",2):f(\\\"\\\"}/****/e3a^15^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"),s[999999],*q=s;int main"));
$write("%s",("()\\\"\\\",2):f(\\\"\\\"{int n,m;for(;*p;)\\\"\\\",2):f(\\\"\\\"{n=(*p-5)%92+(p[1]-5)%92*87;p+=2;if(n>3999)for(m=(*p++-5)%92+6;m--;q++)*q=q[4000-n];else for(;n--;)*q++=*p++;\\\"\\\",2):f(\\\"\\\"}puts(s);return 0;\\\"\\\",2):f(\\\"\\\"}^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"))\\\"\\\",2):f(\\\"\\\"{s+=^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"00g,^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";for(m=1;m<256;m*=2)s+=^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"00g,4,:^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"+(c/m%2>0?^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9)"));
$write("%s",(":f(\\\"\\\"\\\\\\\"\\\"4+^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\":^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")+^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\",^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";f(s);s=^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"4,:,^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";\\\"\\\",2):f(\\\"\\\"}f(s+s);for(c:Base64.getDecoder().decode(^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\""));
$write("%s",("\\\"kaAREREX/I0ALn3n5ef6l/Pz8+fnz58/BOf5/7/hEX/OZzM5mCX/OczmZzBPn5+X/OczMznBL/nM5mZzBPu++fPPOc5zngnnOZzOZgnBMGAW7A==^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"))\\\"\\\",2):f(\\\"\\\"{c=c<0?256+c:c;for(i=0;i++<3;c/=8)f(c%8);f(^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"8*+8*+,^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");\\\"\\\",2):f(\\\"\\\"}f(^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"@^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");^1^\\\"\\\",4):f(\\\"\\\"'|sed -e^1^\\\"\\\",4):f(\\\"\\\"'s/^16^/^32^/g^1^\\\"\\\",4):f(\\\"\\\"' -e^1^\\\"\\\",4):f(\\\"\\\"'s/^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\"));
$write("%s",("\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"/^16^q/g^1^\\\"\\\",4):f(\\\"\\\"' -e^1^\\\"\\\",4):f(\\\"\\\"'s/.*/print ^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^8^nquit/^1^\\\"\\\",4):f(\\\"\\\"'^3^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")\\\"\\\",2):f(\\\"\\\"}^1^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")\\\"\\\",4):f(\\\"\\\"');\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\").split(\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",64):f(\\\"\\\"^\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\"));
$write("%s",("\"\\\"\\\\\\\"\\\");for(int i=1;i<a.length;a[0]+=a[i+1],i+=2)\\\"\\\",2):f(\\\"\\\"{a[0]+=\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",89):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\".repeat(Integer.parseInt(a[i]));\\\"\\\",2):f(\\\"\\\"}System.out.print(a[0]);\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";FORiTO UPBtDO INTn:=ABSt[i];print(REPR(50+n%64)+c+REPR(50+n%8MOD8)+c+REPR(50+nMOD8)+b+\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"J\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"+a)OD\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"while(!=(S:length)0)\\\"\\\",2):f(\\\"\\\"{\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f("));
$write("%s",("\\\"\\\"\\\\\\\"\\\"trans c(S:read)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"D(c:to-integer)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 35 39\\\"\\\",2):f(\\\"\\\"}\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 24 149\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"interp:library\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"afnix-sio\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans o(afnix:sio:OutputTerm)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"o:write B\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");end;\\\"\\\",1):f(\\\"\\\"\\\\\\\"\\\")\\\"\\\",1):f(\\\"\\\"nsys.exit 0'}\\\\\\\"\\\")\\\"\\\",0)]]></xsl:template></xsl:styl"));
$write("%s",("esheet>\\\":s.WriteByte(Asc(c)):Next:End Sub:End Module\")\nput=s\nprint\nqa!"));
end endmodule