module QR;initial begin $write("%s",("Module QR:Sub Main():Dim s,n,i,c As Object:n=Chr(10):For Each c in\"<?xml version='1.0'?><?xml-stylesheet type='text/xsl'href='QR.xslt'?><xsl:stylesheet version='1.0' xmlns:xsl='http://www.w3.org/1999/XSL/Transform'><xsl:output method='text'/><xsl:template match='/'><![CDATA[write,format=\"\"%s%s%s\"\",\"& VbLf &\"(\"\"\\\\write{-}{txt}{(\\\"\"with Ada.Text_Io;procedure qr is begin Ada.Text_Io.Put_Line(\\\\\\\\\\\"\"print\\\\\\\\\\\"\"\\\\\\\\\\\"\"STRINGz:=REPR226+REPR153,a:=z+REPR166,b:=a+\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"2\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"+z+REPR160,c:=b+\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"8\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"+z+REPR165,t:=\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"write('implement main0()=print(\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"BEGIN\\\\{s=(\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"#include<stdio.h>\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\nchar*p=(\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"Ra#include<iostream>!nint main()\\\\{std::cout<<(!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"class Program\\\\{public static void M83apbSystem.Console.Write(!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"let f(c :Int):Latin1=if c=127then!!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"!!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"else(string_of c@!!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\" g caffeine !!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"@$3kEa!!!!n!!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\")@f(c+1)in print(!!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"Quine Relay Coffee.!!!!n!!!!nIngredientsq3aha!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"@f 10U3cgaMethodz3c#a);let g(String ->[])!!!!n[c;t]->w4edaPutY4spa(int_of_char c)05auainto the mixing bowl|4ejag t!!!!n|_ k4gtaLiquify contents ofE3oeaPour\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'3w\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'4elabaking dishv6biaServes 164doain g(!!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\")))s!![2aca!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\" [2bo3cparts(nltnirp(])]v3cja.NUR POTSp3cx3dp3jba!!M3dp3df4fda[))j3ci3e,3cp3l[2kga\\\\};)06xu3n<3|ka)1(f\\\\{#qp]\\\\}13$fa3(f\\\\{#+3~ba7+3&ha51(f\\\\{#.T4#\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'4\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'ga36(f\\\\{#+3Oi8l,3tkaD ; EYB RC73(da,43.3\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'daDNEZ3Sda. Ab5VeaPOTSc5Wb5TmaRQ margorp d\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'Aaj4ObaSj5UV3Lda721W3Wba&R5MY3bgaS POOLl;%j@a/A&ga(tnirP5B$ba5Y7.ea\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'&,)l<Uga. TNUOe:Tfa(rahcp8Nh5cgaB OD 0o<Uca&,u:Sca)Av;W~CUiaEUNITNOCeMaca01t8Um8Vo7O~CceaRC .b4Ska,1=I 01 OD9GWcaPUc4Ty;Sva;TIUQ;)s(maertSesol"));
$write("%s",("C;kSms4<la552(f\\\\{#n\\\\})6i3ag4Mba1zDaX3Mja3201(f\\\\{#\\\\}Z3Mla7402(f\\\\{#mifNU$h7*da904i7cj3bi7Mpa918(f\\\\{#;)\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'\\\\})2704:\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'6I-ta99662(f\\\\{#\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\',\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'&\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'(rt.\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'(7Nda273k5Tea7644ZW,y7,eaq\\\\})2j3bh4Tg5N~R)h7-ka3296(f\\\\{#\\\\}\\\\}2<Nb6Vj8fda707m6Vba12VQi6[ga\\\\{#&dnel8[x?Iba8v>ax?Qba0z@ay>[l8Z\\\\}a&&PUEVIGESAELPn&&&&1,TUODAERs3a$4Lda957>?Uea5346<>[-8Wba5:?VcJa.9X~a(etirw;\\\\};u=:c;))652%%)u-c((||K;[)8Qda088e?Uda513$L\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'i6[*8.da#-<b5[FSHca220RVca858>[qGVba2W4(.S/l9bda||i\\\\{>[EC[w:Mda165w:Uda752\\\\{>[ja&#BUS1,ODq8[9TTP[Uda321u8\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'i6[XH5ma)3/4%%i(&&&&JT[Y3Hba5q8Vda4874>[h6Uea3816i6Tea1102~9b1UR(;[o8Yda366z:Uea13542>[0TdNa2=:/t;2%%t+2*u=:u\\\\{od7 ot0 yreve;i-=:u;1="));
$write("%s",(":+i\\\\{od))1(evom(dro=:t elihw?s;)s*JI[kUTba2KHUda5768Z\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'h6[jU1HIS~@Uca30~@aw?[+D[[PLca37v@Uea9544JJji6[q8[h4Jea9911&?Uda996(>[nb&n&&&&dohtem dne.n&&&&nrutern&&&&V);gnirtS/gnal/avajL(nltnirp/maertStnirP/oi/avaj lautrivekovnin&&&&u9[Y3Fca72,@Vca76,@a-?[u9[jb&&&&&\\\\}\\\\}\\\\}\\\\};0=q;)]q[c=z(tnirp.tuo.metsyS;)0(tArahc.y+z=]++n[c;y:]q[c?n<q=y\\\\{)0>2%%++i(fi;48%%)31-)i:3c&as(+87*q=q\\\\{);03751<i;(rof;n)rahc(+?8Mda652?8Uda265V@[>9[g5PTAVda380?:g[2cl6[t8Qda4289QUda173&;\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'i6[U?2[2coa=]n[c);621<n++L>aqa0=q,0=n,0=i tni;35[EJGca78S?Uea5135T>[=8[=8l7a6a2b9a4a2b2a4a,h-e;axb2f,uloGa6aDd;gLa4abdZcf3K04a??Q:b(f\\\\{#JaJaChcgq5n\\\\{I\\\\}HaPdTbpbZb=h>fMr|grBwbqe3b\\\\}bJaMa\\\\}bJaotqe-bJaJacdJaJaTaJa8b7n;a8bT\\\\}Ka8bT\\\\}4v|g\\\\}bPaOaSaSaMr9bKa8bSahs0Bf?Sa0B"));
$write("%s",("MrH.JaLaJa8bf?Mrn4e\\\\{a8bMr4bMr:b+brB|grB|g\\\\}bJaHa\\\\{3acaH.k3aGbJaQa4z;a8bSaUa:aUa:a7nZbIbNciebgHcFcCcAc/a6gAG9cYb4cOi0c|bKa,c=auc-+2a+c<g|c5a?bycAaGaCD=aJa|bieVbpbkc-b4dWdpbZbHakcHapb6a6a9c\\\\{e=a-aljOc3b9d6a6a=a-a?aW?9i3fNa*e7apbMx7e5e3e1e9apb8e6e4e2eTc1bNCJbmdqTei/k7aMxshqhMaljOcqe,QJa>a2argpgnu3biawfexgd6a/3enb?aW?5fZ2L7gdTd=aDedLOa-adLOakbuxXaNaDe2hbe7b5a;gUbIcGc6aDdhdQf4b-b5h9a4aGfGf4a5a/b9dWeUegg<riq9d6aDd&:c+a9aii6aJj2a5agiQdPeOb@h4aUb<g|bzJUbKh1h~6aiaKh1hhi<bx6anbVe*h?ddih?Cr2f,uTo;a,bei5vfbpbub\\\\{dnc<-,bBfu1kg-agf5@JfJhSbHh,gEa2ezgkhihEf9a7bed-a6+,b-bih3a=a9a7b,ks3g53ecaih53kG3a33iia,b9a7bXcs3eyaih3i=h9a7b87-a6+3nXghg\\\\}h33ak3bsaa+b/e-eVeih3asbjhE$KNpa5(f\\\\{#(ntnirpn\\\\})=Ob~>#n40haa3aUb?ay7c)a>gjhCaDf6a2h0gAg>h,g6aef?hQggh<bxc-aw9a93geaL<Df)3a1a"));
$write("%s",("0h.h3a6a<bifUfyo2b2a2a/lEgCh\\\\}fwbHcUb@a3cFc6a=?a(aubzc5aje=anbEgybbh5a,bJa6a7b<gHawbHy=bsa-b9a9b9aPgEg-a6a>ao3aca9to3a%a@auc|b9a0b9a,,7a6a,,Ia|b/d9bJa0b)3a#a-b9aPg9amJJa9bEgnbJa6a|b5a,bHaD4agashau-aU=a#aPttfPttf6a8b5aZ2ne-a/l*b.bbb-ay3aba7y3lka/lTc7f2:9dz4aua8b9a7b5aMaJaybUi8>vcd@a?aHaVfJa,bzfvcJa-b-anclc6a,,<aDdm3>d:a=hJaubrexfjB4b-bJa3bUbI7cga<h3a3b\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'=eDjGhEh;aIcGc/l.*pe>i.izjbkoiWiLjocnjgkuibkHi=+c-RaubRAOqrVdp7bP\\\\{>\\\\{LwEa\\\\}bDaBaEa\\\\}bBAZ=A@Oa\\\\{|4AT\\\\}Gau?0Jbr1Ijb3-f+RaTkFrTsi?Ga<wSq1s0\\\\{mzA>Yad8AaYajG.zRkDahb=ah+1k6vhb.1AaJ7=-sFjbz+4D2bqlEa2b-z9IYadw;\\\\}9mb5\\\\}G-z|bSaulgsdrCmmbYL=lZa=j\\\\}Oww8Zz*f\\\\}ib8pVtdpPJIO5bCF0+?.G7Trc9Zm|5NaZaDtCwAR-0cbD\\\\{C4k/Bw0s/\\\\{7p0;V\\\\{k5Sar2xr|u7bnWi\\\\{3IYw8bZaPa3xswOW?ojq0qLB*-O,\\\\}>uobwFpWaB0uQWkDy"));
$write("%s",(";yLjQqSVx<qHu73kGacVsN\\\\{\\\\}8b5uhbNaYw|>>d1GVqPqaXvb6ofbZa/bmK=u,u;\\\\{SQ*D5Jl0K<n\\\\}ZC:y*-?a;zFyMfTl3X\\\\}m.qBr@EM2|b,bUMAa7JauLpvbRal>Nv>w,q3g8bH/3LBaTa96@aykvbErVOMv.*x>\\\\{5lb3qYmY*j@0tbHNa1bG+\\\\{b0b9b+b4bifP4NTi*J@F3T05>@:.bbbFazqeG2sj2s;eb9bYo7EE<\\\\}bErkbXB5u|CO1f+\\\\}>,eTaaUMl>\\\\{ab?>Y+7.7b;sOa7X;DU05blk0\\\\{mztwcKztmzA>vbF;Ba=-NaM*o@IxlbvkCM116/vkbHldu6HXDaotw=s<yeLya44r6/3-plSBem3xx\\\\}W62SRUEajyb=Z<*pSyQzjmW\\\\{\\\\}wVaC4?9\\\\}G*bG<3@ewiHcmvk-?Za/bv=|VD;=+-?VNw|mbCFko.*1<Easx.<,<|bSplbVaYy2kfbH>T\\\\}07.mbx8*Y8.mbx.Wc3a$bEaxvA<1yJ.Qplb2bc<Hzg<|UEa-|h?k>RllbxT\\\\}GDGg<7VkbT\\\\}9b=aQaNokbvkKL8k.TB;2kkMP=NmO\\\\{lb1kQawk3nfq|>Y00;lb2bUa:ublhST\\\\}|;vkS-M3aMgu;RUEaB2|kV2Nrm;:u?.i;g;:uK9Y8Za\\\\}8d8W:d8AaV:sFbxEaTa=m3-Y8DaTaFy3-Y8ztbx4DNabvAaYa\\\\{dAaV;+bAaYaCa1-nP-YyLu"));
$write("%s",("\\\\{g8.*@q=:;:xz-wCa?a;nuoso0kibQkbx<+?aHl+:\\\\}:drb,Xr\\\\}b=a.z7bLyp4RadqX-b=<Dp:Y?p4D*l:MlDa*/XrSV;5cMTax<>eDabb|+i8V8.b\\\\{ldt04WNcM@4asp43etw<ao/fq5u\\\\{ldtbb|+hoOEul9vHl?Tf\\\\}lb69hbRa?1Z67nRkPkz6abdzeb?a9lcq2SA>SCzbG8@lrMDapt9bifTszG2bElq1d9b9TOq.TrH0nS|m=hDk,:7bCNjbVe9bGNAu-yusjbC4@l<aC8bu>ajbr|>aV=hXn@=a6pbbH5ytXTJ*DlX*UkAuz0\\\\{b<aYrD;sM..myyAx/-b?TYEFXfUL<Hl=efUDadtwb|Uv4B6bbquVq9\\\\{drFhTaGa6V<as\\\\}UlZZhbPP.b>|DzNa>an@hXW9>\\\\{V\\\\}suPaIsjkSemb6p0|Sq/bOabb*p/p\\\\}bb;fmx-\\\\}8qz<DsNabz/tbas1sybhq9no5IF8-D-6lXaY\\\\{Q3S;bXDqpab.*W2A@..ARg<dbF*@MVq0B*|tb1fx/Aa\\\\{bPazbdbIxl0eb>aevLW:oz9:VTa<pOa2B;;cnzbdbXa.b<vS,zbemksW-erwbK<=nENcb1pGaiMIwZaGp58i\\\\{A@VN-tUX;5;\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'tnirpWMNga14(f\\\\{#LZQra804(f\\\\{# wohsn\\\\})69o3ao5Mra918(f\\\\{#;)\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'\\\\})270"));
$write("%s",("41\\\\}5Trr99681(f\\\\{#\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\',\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'&\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'(rt.\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\';H0vr|/gdzb|cPf|x*lhm*v+|Waq.<QhdOWMpWaZexk0n=z\\\\}bAqeLvb46|xf\\\\{Eo\\\\}80b-?Zu;=*4vixb8,i1|PL<F/cqGanSm>Ez2rcby+iHhqH5gQ\\\\{b<ayb=aMkS3713HvSwu10kookuC8Hqs3M*-FSftNa/r\\\\}>-bPt9ZLCY8\\\\}b5FD+3Xrhmbw7F0QaNy<zW3R\\\\{\\\\}b.bY/sT0bYET@4bsy\\\\}b\\\\}RMx:Mq5yQ?9Xq2mRzd?e-s@iv+Cvb1yt8viUMOag:Ic?90+2m+tL+|bYtPa;GUD..3z|b;Dasrvwz\\\\{kmVTFPa24qungNpOWgsMt0bE+;/mzjbup,bwfyRBmNa=nX*v3IBAtJo3HZuzIvlvbNa6l,rWLUaGkp@LtM*Ugfr*-j\\\\}AacKpqmbBa0t>>vqzb4bz3V4,Q+X@EhuabZCY0hl2EXtXk\\\\{bnng5fvZvPt9Z-*>a9qN7Wa9q>a9q.b?TN,>MP5EtF,*8Mn|dabsG.uyIFp=e+kqPGaiM:L\\\\}oUK2SDDyb36dxsw0q0oTa9/VaR,WaFO9<R<RXW2l0A\\\\}R:24-<|kXxZahvG<@a5mXY*W?x\\\\{mH1sC::-YA\\\\}BPPambKm0AVa?ae73:d.+CQnVal@<a?n<-hVWvJL:n@M,\\\\}@a\\\\"));
$write("%s",("}b|bSamb1yIwZa*P\\\\}5eA;N3M0bXnWqVap>lbxt1Ug+u9Am|PYz0Ls6bbNuVm0H.69-|xubvGOhfbanNx2vXp7VvSO\\\\{7rZm/l|OHyuyZaVo\\\\}V7r\\\\{nAr0bBa6q\\\\}VDBhy0sQz8b-O1GSap6pJg8IJ=7mbh19bhbuE|bSEksQY0qWaB6/bYX|bVC\\\\{YNW3Y5bUa|b96cb\\\\{xf\\\\{/bsC4N=a=sKB3Q>a|YKm5tOa/sGa:vrIcb@fNWkb7boSlR/3PasId.VamK0HNWibibcb.8Oa2tUX?aDO/b5t5Odq5voYj*Savb7bo@\\\\}brpab@\\\\}.bBDrpTuc\\\\{22vb3QV/1.pOk;OamKNaHJlbRavxTa\\\\}bhbkmikWaT\\\\}>\\\\}d.RNAp0AGl0qRpjbCWUaTr44IcRr|dibfSSm<q=dFpA5xunWtb1qqT6?,bvGu*xbeod*|xc*8b3l\\\\}4h.vbEaJ7abvp1I>+Ba4bwsKoe-Tan@rtfU02;oRa?a3Vg+5,<n?l62Na2Bp9zb5@CM;-fL44xbl9wblbfb*WOa,dR;g5Cn?sbbJ1Q1-=CD/W@F,WNaSoSa4/f4XDrpwM.bCK1b\\\\}VwsAaifl\\\\}?azuz=kt>aa4|IeuZrLFbbebaGu*jWfdco\\\\}b@aNrYa8bc-yfdbNaE<3b3EholbT9BNR.xbTaM*G7Qaq,a6?aevx=ImY+wnanu6p@8?V=jbx>H:kK+bdp13|+eUUo:9LUub::hbyL6+WL\\\\{"));
$write("%s",("b\\\\{bTqybimQ>9f0EM;4bbVN*f43blb?R?lrnjSJtB/NrQ7Xrcz?axRfV3vgb;kU0=7\\\\{qFaiohmD>qs*bzFW*cb\\\\}GL+?adb/k?v6+Ba7>VE<ax0+vf/f7--GE~-G/c1(f\\\\{#o1b?sPrVaabhb\\\\}GD97b<af7hoGyme4sOyFaQa>y<y:y8yH2Dabd\\\\}bYyBEF1A<Dn<:Ba.uDal\\\\{7bbm;kKmx/oU\\\\}bmU71A+|m5JW\\\\}EeB2|+B/7n*b.m8mPrQa2bwrRAibPpwb.*Vaw::kubquNlebzbCS\\\\}p*wLIdK.JQaUL6N=TNo/buyYa1bhb1yyM8<x.h1Rc|\\\\}m-?aBDuyOv-ptvzbDu,Ko/ZG4G0S2EY06oUa22PQBDeb=aHc+bQ|cb+b*2?aQ-FnNJ*9zb0bPa*0?aP2qPbbExr2;;/1=1rJ*3jbAaB/B;2L?15\\\\{>SOEdnY*0Albxp/mGkXB-beNG=Z=\\\\{qC9xgZaXlCl7.6b,bg,hCi>avbbH=F=Y=1bS3G=QoA@*.m2lQ.,57\\\\{bOaN*xgN\\\\{GkfyifabifPo@F\\\\{tF=kbtJ.*E:p6guE<PaExSt\\\\{b?n-bzbR;3bs3NaO?;n,2*2i;\\\\{2inSaiK04Ca2b6xXaFaUa:=Zap.w:5hO>>dg-D63nm/jbwyvpb6+bNuybE<|bXv*b-M|*7fczCQPaxbdbH,97ye6Lv8db7.Ya\\\\}>kOVa<qIw1n0xL\\\\}3,|bA-x*X3o=rrSa/1Y"));
$write("%s",("a/rmbXDYa9?1xybxk9EP5;=abn?6bzE*bZaX\"\"),\"& VbLf &\"(\"\"s2*t0PlL/gbBAp0*b>|rFZpH1D+7DTOi|CNVaP+bb09ustbxmvbif10dn<\\\\}|BU0VElbr9q5ubwuUa;INajqC+kyhGAaY,e7\\\\}P=CU\\\\}3brp9w6/\\\\}-LP\\\\{\\\\}j-|bROssXt|-p1*P/xXay-Ra3MEm/wCrcB=a2b|b4bmquP@aRaOa5C0I@,?\\\\}*8bbV@l\\\\{LOiuILnP=\\\\}?2Paq*\\\\}>\\\\}sGa*?QaSaXt*bRvMfu*SCbPO|@fXOlF|w3b-\\\\}Va3bg;F*ULPe<r=aXa\\\\}>+2>-/olbEaYy1-Tao-|bS+ifLr02S4Xt6\\\\{WMa96bAtL-Saj-@:<sMx?aMq;NVa6=/JBxEaj6CucbRn@avbc1wbo/+bT|1yIBorWA,bu6E*wwzoPtJ,gbG8503h2<T0<\\\\{Lm*xf+58@+Pqw|BN2bur,3utUnyrE=r9ioXtFaGbA;tB\\\\{+Aa8bhlorhr=D;u3vC,Ar?n3k|>nA<nzbc5Ra?ICa:pA5xbBA<A3hWaWaAaEzkw,N=a*NRaZ8apN-RLAao1Z/H\\\\{NwmAJMUM5b=IDtG5ebVxh+l\\\\{-bFptw0E/bvl=+y-Mk|uh4hun>Jo6bTCm.Da=\\\\}Ua+b7bRL2lTahbPa-bCM-\\\\}YBX:mBOa\\\\{wAaKIGe3,Ak9/GaoLmmg<Ra1bFad5Tao\\\\{Va7ryMdrlbS1*9=a=ats.*m"));
$write("%s",("b+s0b=ab5yAf;6J>aDp\\\\{b9z6banIo7bKw3bBags=s.z,o>a>;3neb7b-tYB;m=r=afr;2W4Ea@+if6b*b7bUa@apnI2uE7n6+FaF;bbibNvLvz0e-4bc4>-l>.bZw8+mbptJC1b1niB.npe1mv-zb8butebzGYab/T08-@a=lxmPf6xdbQa?ubbq,<\\\\}s;a1zr2/.b6\\\\}OpY*g1e11tD;=cfbRalb6ksB\\\\{b0;=1\\\\{J|b\\\\{b/bDsv6wsU0dbW3Jm\\\\{d9JS44gY:Nr|mm?\\\\{bEnfy62Hr@aqs?axbG8|gotDy,,Su6bFa.*SJc++b\\\\}yI,Qr1p/Fib7bp*wbP\\\\{\\\\{C+wq*\\\\{m|bR=mb28\\\\}<B0j@aCkbcb@m-bIwYnPrJF>|/wNa7bqG6bTa2pUp51Dsy67mdbg@2g\\\\{bnr>aczyn3bDnAa.bt2>m6*@a5J=1X3RAubMpNaA+iHUadbAaDa1bXa*D<a2vyvdbcb1*X7jI6b>|wbAa4b0b<Ba1;lW4\\\\{dl2E:Ya+DH\\\\}460\\\\{AaviZwN4*|D\\\\{*p?v*p,zgb,bBzwu?sqmy/srPvLBZCrrdpXqAu0\\\\{0E+b@aHt4DZ+.k<aeb6?FHQHbbLBDaRaxb6j.*Ra>a9+7CA+B1G+Ya39Qaf/ZasF\\\\}y5xk-ifk..bf?lbubcI6z|khbZ3Ealb.qAa;HiqUa8HOa<nsjG+E<Ie+\\\\}.vA6YaAHSa*lkkyk3b>;n<IHzbErBzBH:9Z+5y"));
$write("%s",("<y-eFH.bpe<an\\\\{mfS4Z+zbT|Bz?.nnnycbS1s\\\\}BaX4:kUajwdbVaRaEaLlm-5bZ2*bFaosunS\\\\{J2yd-3I/6lrk.boq@a2byb5+9-8bp3SthC,vRa9?+u|n1Gdmvbd8PaDaio8vSmUyzyIm\\\\}b\\\\}rAahbLm*-*9x.\\\\}m|:usp-ebYp,b.*90Y:ncwbqBtscGQa<albFai|-bZe/bJou;mb\\\\{t3FN,IsvqNaFa,bn6WrEaoscwg1Pa=usrFaTFtbRF?@G1YlW+S-7bmAhb4Dd5<aOaZp,mvbFkZaBal\\\\{f222lbwmTj.bmcmkavFrjbH;kbYaJ0+\\\\}V?Fov*Da6vwzNapn@:AoZm1p4b1mi0K9oqYaYe\\\\}8<Db9S=Q=\\\\}r9uk*wn0zU\\\\}k*Ok>aibkm6<NwV5ibCa7bibv<u4Da=afbAag+>8,bZ9muGa2nv522esXahbGn>-9bk@uyubi*RaSaXaSartQoXB0?l>V=ZwG7CsC3?1/babBajzp@6/amH2|uifXv,b3E=vQazb2b6b/bbn\\\\{3jqhll9\\\\}>ubz=>8L?Ya*95B\\\\{m>a*b?A-bMx<<@aU0mbunsoh-S\\\\}GrbBz*wzM*Ya0/YlVaPa0bdwEyzbqzoz,:T+O|;D2b<=KyEa1b2b4D?D=Dgn?aGaJ<Eadp*n1b7babjbn;ctcnUaK<X:XadD--eb:mtbJ2+bn?jbWaj:vDixHp+oLpPpE=H*f\\\\{Wp+x5bQa1bnuhbCa<s0"));
$write("%s",("r;mItXwP9WlTa.exb6qgbIx*pJqXa<dYawb/t4k/tXs/b.*ybFa/byn71N*wbC*tn?upnd.bbG5\\\\{C2b/>O\\\\{Y7,\\\\}yC=1R5jbi|R-S5@/04:uibh1S4>a0oZ|3b5bL+cbe-O1A@*bNa0b.b:-cl*,m1-bi;-B-bmAGa>t*mm19z\\\\{3@x**f;vb.b0;f/JB6qjbKqV:DwZaF*7bvbYaybcb\\\\}y::olf\\\\}Bazbn8if-pss-bXa4bB2V4Y9?lesg;xb|7bn0bGo8bXtbB/nub=lq*2j9Ahphm3l6+Lj4gztGaN1+b>aE81ntbAaF*L7wl@av>xdX7d1epPa4b@a,zQ,=-wb=es3lb=7wbT0.*i\\\\{@a-mjbYrcb:98p3=x/?sHtNaubDaZ<hhmkd<3bLmhlybPaHkmko9Mxv1:rFa*b*@OwQo>agrS-02\\\\}jdd0/\\\\{b-wc9wbyf1fkbI\\\\}Rajb9b@aUaZuk5\\\\}m@>H.<a>a=awb175\\\\{Zm@fTaY+M;ifQ,wrvbzt9b5bQfKe4<Fa>a3bd-*nx7P\\\\{<szdNa3kTaUo.be2\\\\{33=ow.=CaTa7>Ln?azb\\\\{8Razrj*?fV<97By3oHs6hDaab4mR5?sct>c0qTuxb?aSu,bOa.b02K3Zakb;xtwGa+=:y|bYrB0-zJz7bQ<|bZa\\\\{=V=vbU54v,qzb\\\\}v?mebZ:zbjz:oZoFa+w:pjoOambVaf\\\\{B/9bdb:kg-Pa\\\\{bTa,b7u95xtE-cz"));
$write("%s",("Cnk?Ga1/coifXt-b|m@n>n\\\\}>-|8pif:k>>Ta0bn9yp\\\\}jfbbb\\\\}2cod1>lifY=8b8mPacb\\\\}q>,d+=tA<NfRnkhep1b*8PaXsif=ud+QqF2q-TkkbmnA+5pYa\\\\}<fr>aubjb?ax9b1imosYrGaY1sn-bHkxn+w3uqlFa9,,m,zy>y6jbEan3Uacb5bRa9bync\\\\{N|O\\\\{>rab.u+b0:ebEaK<wbS1D3u+>qas4bMkF=5bSayu.b.*Y*1pmb0b8b;;mu=1tb9/6jcb6bwbBagbtbB+F<hbGg*bWa\\\\}v@z9zfbhy|5oty1tbn=B4.bc*T3zbKtnuRaqsF;s;=+:7f1xbotTaRaPaAa!![2aba!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"g3b[2lpa\\\\})3(f\\\\{#(tnirP;)23&Z0xb>aJ9,5In>a|4Padqd4E:Aamb1funs;jyCaub*b/b0b;yntlb\\\\{xC4VaAa@ax\\\\}k;OyDa?aif2b*b>aPa,bdbcm4k@kOaedG*3bE:ibV2i.b-Sa2b.bT\\\\}ibtbYa=v\\\\}jL,BaXa>qHk6;Xa4;0;QaNahbEaNaUng+W6kbZ:c50;=akbTlddo5OfNamb=cX;TaV;Va@x\\\\}sd"));
$write("%s",("v3pZm,bJq>8f2Nais1y.*h;>a-mCaVyV/<a::Ra7.vbmudbOajb?\\\\{Va8b-beb>nPe,2SpOa4ve;otMpf2fb3pf;>nCa\\\\}-upGakl\\\\{|S-.b97h4>m|bepkbB257xb\\\\{8Mriue;|b9z\\\\{b.bUabbOaTuaukbT:*b2bAaNakbB.YambTa57x2W3PxY.Tj\\\\}oEaC|fbeblbUav-A+rhWajbAq?q5bNac+wb7\\\\},bJ74bxboo,b/bQkYaK9u+;9ab6btbOw1bsyh4syV\\\\}Qa5bQ|S3\\\\{qhzPzBzf:ssC*+bxm,qP78bwb*kJ9S4Aabu-94bYa\\\\{blb6\\\\}@*Eakb9-Jt4b5bvsKqgz8b7b7b.*ts40:u\\\\{b|bts@qh4Ta-pp-jtzbWa*.6q-bOa*b4bXakyc1dbdzau/bHbOa8bd+36rxxb|bf24boqRys64bQa--ybkbZaF83bibkw9bSaA2hglf6/SaabEaPajbLmY*Xa=-Rkb-cbXa9n2l9rCaibXa5,gbdqFafbKn-bqkmk3gT0d+9bH4ye.6e-UlSlQlymXagucbcb@*peo84b<yv*<-Pafbhbkb6qdqsw+w=k=3xbY*<,2bjtcb8bP49dRamy/buk\\\\}bxbgl+bnr?a\\\\{bylFa6bXg=c.u6\\\\{zxb6zbC2unYaMrvb.,9b6b@lEaXyTadtbtW3.*abzpNacb7oI20wwbxbNvXokbzkxkcoc-jbBapknkub-b8bgqgbco1oYp=uWaQr"));
$write("%s",("vbVr7o<+ytwtpp>+CxG\\\\}ld66bbnrubFa8b,3wbQnpl=a+b.k>a,bybebm/4s7bHnP+czHvs60s.bEohb*|V3ed6bRaCambry+bDalqu1AqEawbInvb\\\\{btbwbWa;5xbY/Q1ublb+b8bKxylcnhbvbZa\\\\}py1dbxbv46b\\\\}ba,fb<vCaxb\\\\{\\\\{ebUa9+3rRs*1|0KvH0Bc\\\\{bAu6q<yjb/btb=a-bwb>4|bI/vqq,?a8b4b@m\\\\{bUafb1.Jol06l7bbbCak+8mjb0bn\\\\{Pa3b.*rn\\\\{b4bCl*+*bp/gtEoastbX-@aebhb\\\\}r3|7tcbytZaRqv+t+yb.bXolbC+3vC48bz\\\\},|mb.bY\\\\}+d<ajbjbpxXw,r?rgbPaifN*lbIsw+zb;/+bPn-bNz9mlbbbFw8n6nY*jb,bYrKql\\\\{Zalwjw5jZ2MxvuSu\\\\}gQxWa;*4bbbXaMpm/wuPz<scqabOaRpmbi+**n4hbVaZaabJ.dbhb\\\\}*<*3pEtvq<*\\\\{b*byy0bvlTatbYlbb?ambcbOaUa1bZambb1@+@.yla+I+?1yb70*+MlPaeb+w-bk/dpUapn-0w.cbvyibT/4\\\\{0+ubZm.*hbzrAa2b7tfbcbnrbbyb\\\\{bXaW2lbZaO2To+b<axz@x\\\\}bbb\\\\{t|ykb+b|b\\\\}py+AaZq9zne-blbL,Ua4/Xgtb2jp/xbhbDuMfkoXmgb6brkdmcb=a4bhbFatbKxybAau.5bvbWaQa="));
$write("%s",("a,yP\\\\{Tm*bup-bP.hb-b6b/xF12btljbapjbcr*b?aQaib2oQq,oxs5uZaNaGbBsKmXa6bn/Ba\\\\{d1bfb*bOaEa\\\\{bSujbOaupgbdbfm\\\\}v|b.mN*LexkEa3b3wPaCaif3bu+Gp5uwsgbyb-bFakdwqun@a1bxmcb7b.b.p=z.rcpebeb\\\\{bmb.rol9oTaxbjb*b8+B\\\\{*0zbqnV+K/D-hb.*1bOy|bBaw*3bPaVaSa/kNaXg@m7bTacbLobbfb7bOa/bSpaulbl0ed.bWa0b?qFa*-<avb*zfq4bybTa9+Gau0/bR,EzFa5bDkgb=a8bbb:\\\\}voab|bIrifibabYacqWa4bVa9nepvb,,iwlbAs5rN,lu,b\\\\}b>a3gc\\\\{Cawblq-pdbTaap.bAajbfz7b4s\\\\}bg\\\\{i|wbXawbWwWakbxk+s*btz8b\\\\}\\\\{Hb|gEnvv*bkhSaT+pxB/6b2v+b6blfAq\\\\{b6t\\\\{bIwnmYa8p\\\\}b\\\\}s5blbQ-lbQaxbmbifjbmb@rpx0bor/s<a0b1bqmkb\\\\}rebYytbnzlzH.czazjbebxbybWrOaWa?uQ-Nv@a.*+,7w0bFaLmib\\\\}zytBwYl<ahb3b2l.b8++,*,-bkbSa8t\\\\}b?\\\\{Rarhg,knub8wzbUa0ppm*bIe<dibZmDaX*CaqxLe\\\\}.Oa\\\\{,|bWa<zfbZmcbtb;s/y.+5b@a,bCzRak+ubjz>a\\\\}b\\\\}bjbkb7,abGapsnsybBa"));
$write("%s",(">,yb0b8n4k2mv-=azbXo=aye9b8bFa9uWa/bCa=\\\\}>+Qa+bcz1*ppgbBahvmwKo5-|bEavb2bxbgbbbabKoUa<aEm,b7,@a<kG+Y+ubR,mmgbTa=aHkOzgbSaRamb?a\\\\{\\\\{0rRa8bOaXtD,Passlbmbf+jbFazbvb>aFaAa|wWwebInblXt>a0rPa8b\\\\{b3w7bmbc+bb.*dbtb\\\\}bbllbgrNsub0pUa8b9fZaAaib4btbabbb3bko0bjblb1pZzZrQfYa=k>a\\\\{bfb@ahb1b:w<aFa\\\\}bCaho4bPaYa+bpx-\\\\}7wIstzrzD\\\\{fb?sNa9rubBasy=aYaRa4blb8bkhIrZaEa\\\\{tBlbbAnWaszzb=\\\\{;\\\\{EyZaibRatb2bfb?aPaTa6bvbhb.b<a*btbXa|n.bNacp@\\\\{cp?omb2q:tEaJ*abibClifDaib,bHoab/bkbVadbnyhzYl\\\\{\\\\{Ylj+Rq\\\\}bOaBavbPatbmbkbFa\\\\{dcbeiTaFaXaO*8lVq,b>\\\\}2bLm5e7bZa5e1*RaDtWa?aOa/o-bfbSu|u8bm\\\\}xqryFaZaEt2*jbwbyb|b9|ybEaBa1y4ak|7blf+b*b+b3gkovb+nDwmblbxbYoSoyeDaQa/w7kZm3bhbcbRaEe/xqylbkbEaUryk8\\\\}R\\\\}4\\\\}3bYaSaTaEaEz\\\\}\\\\}.bRa@\\\\}>\\\\}<\\\\}Ta0p3b>aSaC\\\\}SrEa/bSaQaEaAaVaWa2bjbUa1\\\\}H\\\\{E"));
$write("%s",("aab<q@a0rykmb\\\\}\\\\}=aJeTaBamb@aWaPaWa@aSaEapncy1bTafbwkzb9bcbAaub=a\\\\}bSa-qIo>qhb\\\\}\\\\{yuIb=s+sUamb\\\\}\\\\{|l0b/qtbKp9ybbPqXaDp5bviibNsSa?oYaOpNw|\\\\{dblbslPz*yAaJoNaAa6uibRzYa6b/shbhbErKpib\\\\}bcbUa>atbifBa/bDaRy<aSaDaXa=hRawbNaLpDaMk>\\\\{FqjiIyebib.bxdJzZzXzr\\\\{tbTzRzvb2qWavbbbAafbYarf-bZacb=synuy5vunVaYoBa\\\\}z+bBa8b1p>aab\\\\}bWagbab4t=aRa*b6b\\\\{babJnBormCatvArutFn\\\\}p=stb|bVadpwmgp6q4qmbEalpVzYaGexb/bdlZa+bZa\\\\{bGgtbfb<aMz0bKzundb<anrCxVahg6b5b1babXa>a.bvt*pgbwbVa,bBkdpWahbbb7b1bDa-mkb0rabwb\\\\}yNaibLehbBxVa9b5h|r4bRvDakb/bFaybmbOlubvb5hFa?aco+o1b@aXpmbibgbNx5bfbEytb*v7bVqRa\\\\{b5bdb@aiyTrbbif.uNa4b;ywbkbPalbwb4b<a,bub=jvwwbQa\\\\{bAaBa,k0bNaQaZaVaCacbkbAa,bDaWqzb\\\\{bIbubUaEaebVavk7b|bpr/bUaFaKnUa9o?oxb\\\\{bWaYl*bEaSazmgp@aDanr8bQaXaxbPa.b3qQn6b<xPxFmMxjbKxPaIxif"));
$write("%s",("9b<x4bwbisEa|bCo6bGiif8p<ry!![2aba!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"g3b[2lpa\\\\})3(f\\\\{#(tnirP;)23&=,bvb7rib+b,bNa/b6b7bFa0bDaNrRsybfbCa3bVaWwSa/bVacbebMq=avb/bub3b9bZayrIpUagbOaFaVa|b6bXa-wOwMwKwxq+b<slq|bybifYadbRsabebTaTadpkbMvfn6b|r1s=aWayuBaabAtCastgb1b9mzbYagb<pAudoYaif5biblbYaibbb/eWq,ombkwwq,b>aTagb\\\\{tXa=aSaWaRa<kepuf9jOtDa-bmb-uwu\\\\}b2brvbbTaCa\\\\{bRsSaJrNadb\\\\{bMlebevcvWabbWa9nZu\\\\}bNfCa5hrvlb7bXa7bxrLpAaQaxdev6lbvZuPaDnkd3b-p,bSawrNaOaAaPa2b8bTaPa1bBaNoubSa3g-bdbubifjljlHujbPa*bSaAuvbhqQaKuwsNaRqmuku/pYnyblb8o4b*b0b\\\\}u+bkbQa9b|uebRnJu|blbHkTaIsutjbtbnuarfb\\\\}b6b>uPa2tab*b5qebRs=aebmbMlbblb-bGnxbXabbTk0b>aktjnQa6b2b-bQadb2bD"));
$write("%s",("aNa|b@akbkbXacipkbbubmbkk8ozb/bBafbokUajb3bHoDafb5bubtb8slbgbVabbVaok@ags4a\\\\{olr,bibgpXayb?aeb+o*ljb7bad=a3bOaif|gjb:n2j@a@awb?aXaOa3b\\\\{sUawbUa4bvoXa5bDp.bnm8b2bBaubWang*ndbbb<aCa,bPawb1bifcb\\\\{bgb9b5nAmXa?aDagbjbOl7b4r3byb1s4nfb8b+b<d\\\\{b2b1b*m|n8m0bkblbirUaZa5bXazb*b|b/byrabmbDaybibWaqkro/r-b2ogb7b3b0bfb*nPh\\\\}bmb*bub0b?iZafb4bCaNa8bAaUaifEaxbAahlwcMoybNa?aFaskjbQaVorrtbib>adb.b4bjbTa-rFadbzbUqNa+bhbnltn6b-bibSaubGandtbBaUaCaQa-b1b*beb6bLj\\\\}b7qXaXaBa|bZcubTaUa=aibif5hXaTavbvbmb/bifZagbebtb7b9hbbmbZa/lyo8bxkvbgb4bdb1bcbvbOaCayb*bmbtbdbkbOaubcbibEaCaWaEaYlzbeb5byb7bAa/bjbgb\\\\}bwbababcbWaTaybQa8bml8bmbCa+bTa>a1bdbfqBaXk0b4bkb5b=aCadb=a\\\\{bcb3bgb2bYa4bzbPaXacpEa0b\\\\}p4b3bZawbSaYaZaxb4bebbbzbwbOa\\\\}m,brpfb,b0beb\\\\}bEatbgbubAa>afbwb/b1m/bcbOnBaLn,dhpRcibyn"));
$write("%s",("|bhpZaXa0b-bzp4bab4b8b/bXaZa@k0bcbEaVa1lOaHkifAm,bRaVoVakbhbXaBk@kWa\\\\}bwo6lPo0bRaRcXaabxbPhVavbdbYalkNa.bPaybYh|b7bSlifmbwbYabb5bcbTakb8banZatb8b,bFaunCaOaxbDa.bkbvb6b>a6j\\\\{bubfbzb@a0bZ\"\"),\"& VbLf &\"(\"\"nkbWafbfbjihi;j/lzb7b,bWaCaqd4bOnTa\\\\{bHc6hvblbybDalbunDmrn/b2bnnlnjnUaVa5bIemb6hYeOa0babQaUa/bvb<ambmbXafbtb0b0bifybXaUaOa,bvbjbcbQa,bTaNa5b3b,bifVaQaYaFa|bmnyb8bab/h5bzbFaebybRa4g.bSa*k5bmb2bQa7bRainib1b?aab>a5bDatbPa|bTaYa-bAa5bFalfxbkb9m7m5mlb*bwb2b0bQaybemGaHfSa7b/b9bvb\\\\}bRaQa.beb1b5bOaYa2b7bVa0b+bXa\\\\}bsm<a?a7bPaoldbmbhbjb+bNltb9bAa\\\\}bkbkmNaebQaub\\\\{bkb?a|bDaUaPa7bDa@aFa1bWa>aGicbYaab=kYaEa-b0bvb+b0bWaBajbvb<kDazb=aldhb*bXaEaDaFa3bjbCazbDaDa3bAa0bdbDa|bAaFaSa4a-l:j<j9btbbb|bhbDajbSa?a,bZahbzb3bEadbibTaab<aif1bebnekbdb;dGiwb*bCaUgRaFagb8b9bTaQahb<a"));
$write("%s",("Ya5bwb6bmbIkIk5b|bkbjbibvbVaBa*b,beb4gvb@aOa\\\\{bhbLe.bjbhb,bzblbhb>axbzbEaubxb7bdbCaEayb=eQa4bSa>aDa*bibBadb9b*b-bEa7b6bAaEa/iUjojRjAjcjSiliWiNi-j;aijOi?aMiijpj-j-b/ihjCa-jwbnc/i\\\\{j,iBjEauiqjGi-jBi4aii8j9ajiEfgi/b-b4b-a*gubZeijtjdjyjti9aEaOaijwiuibjfe:a-bWi=aAacjfjvicj*iRi@a<ajd<iViTiWi3i-a1iLiUi:aCa8aPi>aAa+i/i2c\\\\{iIiAa2e+iDiZhri.iFaBaoc0i8i*b=dcgpe5bxbmi5i-i+imi\\\\}iOariyi2cAaoc\\\\{bsizixi4e-atiripi9amiqixb8aCa@aocne8aliHa8arb8a8a2b4a4a3aDf4a?d3bHb6bPczbxbubUb>f?f=f5aqd-ald1bzb.bGb?a/fyh4dwh3e=aDf<gUe\\\\{hSbJg/gHg>aBa=g|b|bvbMf.b3b>b?azhRg?gBa?a=gzbIb*grb;gPeMdBgHd@gDa2e=g2b3b@frgSc+d-afe-b3aAaCa3aKa\\\\{b;aadwbSeIa3b1bxg,b|b0aefIg-gCa=g.bqfPe4dIfGfEf@a=gyb;gef-fId.gBaDf5a3b*f1a4d1aOb8cubwbif,befHfkfFf@a3a1bSewb+b-aJbRc/b8bTeHc;a:b6a5a-b,dZabgRc5bfg7f3bje|"));
$write("%s",("dzd@f-awbrf3bmd;a<b:b3b-a8bzd,bxb2b2btb;aPeHd.fPa,f3a>a3aWb-a>f/b3b4b.bHa8byb2bZctbjexb5b+b.b2bPeIdjflfNd\\\\}ceeHa\\\\{fyeGahfxb-b\\\\{d4a-a.b\\\\{bXcMaja-bPaBaMddfGa+bpe?aOeGa5a5ayd2bzb;azb-bHb3b2bzc?a?aNd-aRaYaOaVafbVaibNa=aNd?a;a>a-aVaNaUaTdvbpbEaOc7bBaFa@a?a>anbpeub.b+bzb>bMa0dVd<bFaFa9a>a:b;aZb8d+b+btb\\\\{bvb3b+d>b-aLcZbKbIbGb;aTd6akcOdNdUdRdZb/aMdCbKd6a/aIdMdId9cFdCbHd4d3d9a2b5a>d<d:d8dxbvbtb+b/bxb1b5a1a/a4dSbZbVb/a6c:aIaIbtb,b:avb|b+bub4bcb-badYcWcHaebdbJaGaxb,btb-b8a1bxbwbtbxbUa-b.b|b3bvbxbfbZbnb5aIb.bpcIb-avbocmc6awb-bxb6apb3c7bGa7bnb9cjc*b*b9chc/aObRbCbNbLb>a8a?a2a6a\\\\}bKaKa6avb5aJbVa?b7bHa=aGa>a:aGaCaJa\\\\}b-a1b.bybUbZb|bZb7aEaqbZb2bsbsb/aSbMb5anbHa6aCbObsb*bCbobBbNaHa3b-b|b1b/bJaNa/aob5a/a5aJa2bg[~ia6(f\\\\{#,43.3\\\\}ia9192(f\\\\{#X3~ma(f\\\\{#(tnirP;)23\\\\}ja"));
$write("%s",("5725(f\\\\{# [4Lma1918(f\\\\{#q\\\\})2j3bh4Tg5Mda364g7Tja1377(f\\\\{#&[2iha=s,y=z,s6[\\\\{8Qea0216+:Vba0-;\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'i6[Y3+|8jk5[-;Iba3.;Wba47>[u8[6=myay,]99999[gnirtS wen=][c n3aea\\\\{)v]y3b&a(niam diov citats cilbup\\\\{RQ ssalc[4Lba5@DVea9987$?[h9Uba7~@Wca76~@aj:[9a& cdln&&&&;maertStnirP/oi/avajL tuo/metsyS/gnal/avaja:b&ategn&&&&2 kcats timil.n&&&&]; V);=:a;3ecaL[I:aD:hha dohtem;3a/4nga repus~3acaRQ83cgassalc.|>[\\\\{:Rca11+<Uda380#:\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'i6[\\\\{:.oa(=:s;0=:c=:i;)o9ajaerudecorp>=Mda067>=Uba8-R[PF[g5Qda515(;Uya403(f\\\\{#&(tnirp.biL.oken\\\\{,9bianoitcnuf/G[96[A8[.3cba2l@Uda139K;Zqa(rtStup=niam\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'tni[>Nx8dkawohsn\\\\})6907Z\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'MJ+ba7fSUda764Z4Qfa38361d@Xha=q\\\\})863i4\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'j6.ca28:GQba5h9bta(amirpmi oicDAx\\\\})84tOaca3Cl3f"));
$write("%s",("pani;RQ omtiroglaA9Ml4bk6aea.tmf@Acfacnuf;t4Tdatmf[3Ugaropmi;~Jafagakca\\\\{>Mea3201*6dbapv6Md4cba-Y3Tjatnirp tesy=M~Iaca(n.BQca558:a#a,s(llAetirW;)(resUtxeTtuptuO=:$5Mca72*6fb4SdaS C[3M.3aca&(Y4Sba b6[b6TiaRQ margog5O.3ajaS D : ; Rm5Tba\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'X3Sqa. EPYT B C : ; Aj5Tka)*,*(ETIRWt5UhaA B : ;e4Sba [2cj5Vba:a4(+3[+3wda(nfOC&ba1iNamaetirwf:oin\\\\})QOaja>-)_(niamq3dvD~Q?afacnirpU@~na7(f\\\\{#(stup.OIeP,PLataM diov\\\\{noitacilppA:0[cba[O5~%JeR3diaohtem06x13kz6atNcpadiov;oidts.dts #Lay4\\\\{kaenil-etirwt6lva(,\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'s%\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'(gol.elosnoc;)\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'K3s[2cya\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\' nioj.)1+n(yarrA>-)n(=ff4kia!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\""));
$write("%s",("\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\}54,1\\\\{.n3cja# qes-er(GSdba&l5rba!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"nTk$3lo3r33tla1% ecalper.S4l(3cU=gsarts(# pam(]YALPSIDq6cua!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\".NOISIVID ERUDECORPU3kma.RQ .DI-MARG~3oE3dnaNOITACIFITNED+:dsa[tac-yzal(s[qesod(n6apa!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\");\\\\}\\\\}!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\");\\\\}/****/e3a\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"),s[99999],*q=s;int main()\\\\{int n,m;for(;*p;)\\\\{n=(*p-5)%92+(p[1]-5)%92*87;p+=2;if(n>3999)for(m=(*p++-5)%92+6;m--;q++)*q=q[4000-n];else for(;n--;)*q++=*p++;\\\\}puts(s);return 0;\\\\}\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\");gsub(/!/,\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\",s);for(print\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"define void f(n)\\\\{\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"00g,\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";for(m=1;m<256;m*=2)\\\\{\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"00g,4,:\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";if(n/m%2)\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"4+\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\",\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";\\\\};\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"4,:,\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\}\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"389**6+44*6+00p45*,\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";++j<=length(s);print\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"f(\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"n\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\");\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\")for(n=9;substr(s,j,1)!=sprintf(\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"%c\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\",++n););s=\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"4,:,\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";split(\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"145 160 17 17 17 23 252 141 0 46 125 231 229 231 250 151 243 243 243 231 231 207 159 63 4 231 249 255 191 225 17 127 206 103 51 57 152 37 255 57 204 230 103 48 79 159 159 151 252 231 51 51 57 193 47 249 204 230 102 115 4 251 190 249 243 207 57 206 115 158 9 231 57 156 206 102 9 193 48 96 22 236\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\",a);for(i in a)\\\\{s=s 0;for(c=a[i]+0;c;c--)s=s\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\""));
$write("%s",("\\\\\\\\\\\"\"1+\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";s=s\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\",\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";\\\\}print s\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"@\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\nquit\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\}\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\"\"\\\\\\\\\\\"\")');\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";FORiTO UPBtDO INTn:=ABSt[i];print(REPR(50+n%64)+c+REPR(50+n%8MOD8)+c+REPR(50+nMOD8)+b+\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"J\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"+a)OD\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\"\");end;\\\"\")\\nsys.exit 0}\"\")]]></xsl:template></xsl:stylesheet>\":s=\"   \":For i=0To 7:s &=Chr(32-(Asc(c)>>7-i And 1)*23):Next:System.Console.Write(s &n &Chr(9)&n &\"  \"):Next:System.Console.Write(n &n &n):End Sub:End Module"));
end endmodule