module QR;initial begin $write("%s",("let s=(\"Module QR:Sub Main():Dim c,n,s As Object=System.Console.OpenStandardOutput(),t()As Short={26,34,86,127,148,158,200}:For Each c in\\\"BasmCBBBCRE`F<<<<C<`C<B`BBD#CXwasi_snapshot_preview1Jfd_writeBBEEDCDGECB@IUDHmemoryDBH_startBDL|DRBAC BAJlACA4RB9MiCD<AERCA>D!BE@ABRCABRCABRCAJ!CE@ B-BB CACk:CvACqRC COBMADRCACRCADRCABRCABRC BACj:B-BBOBMADRCADRCADRCAFRCMM}CBABM~(BBBCBBB,BBBDBBB0BBBDBBB4BBB=BBB?BBB;BBB ...\\\\t..\\\\n..(module(import :wasi_snapshot_preview1: :fd_write: (func(param i32 i32 i32 i32)(result i32)))(memory(export :memory:)(data :\\\\08\\\\00\\\\00\\\\00$:))(func(export :_start:)i32.const 1 i32.const 0 i32.const 1 i32.const 0 call 0 drop))\\\":c=Asc(c):If c=36:For c=0To 11:s.WriteByte(If(c Mod 3,Asc(629795.ToString(\\\"x8\\\")(1Xor 7-c*2\\\\3)),92)):Next:Else:n="));
$write("%s",("(c>124)*(8*c-40656):Do While n>127:s.WriteByte(128+(127And n)):n\\\\=128:Loop:s.WriteByte(If(c<125,If((c-1)\\\\7-8,c+66*(c>65And c<91),t(c-57)),n)):End If:Next:For Each c in\\\"<?xml version='1.0'?><?xml-stylesheet type='text/xsl'href='QR.xslt'?><xsl:stylesheet version='1.0' xmlns:xsl='http://www.w3.org/1999/XSL/Transform'><xsl:output method='text'/><xsl:template match='/'><![CDATA[sub f(s$,n)print(s$);:for i=1to n print(\\\"\\\"\\\\\\\\\\\"\\\");:next:end sub:f(\\\"\\\"write,format=\\\\\\\"\\\"%s%s%s%s\\\\\\\"\\\",\\\\n(\\\\\\\"\\\"\\\"\\\",2):f(\\\"\\\"write{-}{txt}{echo -E $'(\\\"\\\",1):f(\\\"\\\"\\\\\\\"\\\"with Ada.Text_Io;procedure qr is begin Ada.Text_Io.Put(\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans B(Buffer)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans O(n)\\\"\\\",2):f(\\\"\\\"{\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&"));
$write("%s",("Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"B:add(Byte(+ 128 n))\\\"\\\",2):f(\\\"\\\"}\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans f(v n)\\\"\\\",2):f(\\\"\\\"{\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"O(+(/ n 64)107)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"O(n:mod 64)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"O v\\\"\\\",2):f(\\\"\\\"}\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans D(n)\\\"\\\",2):f(\\\"\\\"{if(< n 4)\\\"\\\",2):f(\\\"\\\"{f(+(* 6 n)9)48\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{if(n:odd-p)\\\"\\\",2):f(\\\"\\\"{D(- n 3)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 27 48\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\","));
$write("%s",("4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 36 11\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{D(/ n 2)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 21 48\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 48 20\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans S(Buffer\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"STRINGz:=REPR226+REPR153,a:=z+REPR166,b:=a+\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"2\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"+z+REPR160,c:=b+\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"8\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"+z+REPR165,t:=\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"class QR\\\"\\\",2):f(\\\"\\\"{public static void main(String[]a)\\\"\\\",2):f(\\\"\\"));
$write("%s",("\"{a=(\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"write(\\\"\\\",4):f(\\\"\\\"'implement main0()=print(^1^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"BEGIN\\\"\\\",2):f(\\\"\\\"{print(^3^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"echo ^1^\\\"\\\",4):f(\\\"\\\"'f(s)\\\"\\\",2):f(\\\"\\\"{System.out.print(s);\\\"\\\",2):f(\\\"\\\"}s=^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"389**6+44*6+00p45*,^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";for(c:(^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"#include<stdio.h>^8^nchar*p=(^15^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\""));
$write("%s",("\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"Ra#include<iostream>^16^nint main()\\\"\\\",2):f(\\\"\\\"{std::cout<<(^31^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"class Program\\\"\\\",2):f(\\\"\\\"{public static void M83abbSystem.Console.Write(^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"Quine Relay Coffee.^64^n^64^nIngredients.^64^n^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");for(int i=9;i++<126;)[3pva$^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",2):f(\\\"\\\"{i\\\"\\\",2):f(\\\"\\\"} g caffeine \\\"\\\",2):f(\\\"\\\"{i\\\"\\\",2):f(\\\"\\\"}I3b54rja^64^nMethodv4f#aeach(char c in(^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\""));
$write("%s",("\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")))^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^32^[2al3dp3c[2cs3c,3l[2k@3kqa^31^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")s rts(ecalper.h3eja^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"     53c4a SUTATS(egassem^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"rts(nltnirp(])]^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\".NUR POTSu4cba.C3dh3dX3bba[65bX4df5lp3lna\\\"\\\",2):f(\\\"\\\"})1(f\\\"\\\",2):f(\\\"\\\"{#\\\"\\\",2):f(\\\"\\\"};)06xt3dba;+3nna3(f\\\"\\\",2):f(\\\""));
$write("%s",("\\\"{#qp]^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'[p]#3sv3r23)ga7(f\\\"\\\",2):f(\\\"\\\"{#.33)ca51h4-ba1S4w23F?7d33&r7u53sda,4353.ma^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"' D ; EYB RC"));
$write("%s",("L4/v4+ja36(f\\\"\\\",2):f(\\\"\\\"{#DNEm4[m4ada. A~5[p4deaPOTSn4[#5e~5[o4boaRQ margorp dnex4[x4abaS*5[m4c2<[ca91j4[j4eba&%6[l4bgaS POOL)<[:7dba^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'j4[j4[j4gda&,)(6[?>cga. TNUO<7[s4bfa(rahcg:[(5dgaB OD 0B>[t4cca&,,<[,<aca)A36[;=e6=[.6cqaEUNITNOC      01z4[c9c,5[W8dK7[aGeeaRC .p4[p4aka,1=I 01 ODt4[TKecaPUq4[/I[6<hva;TIUQ;)s(maertSesolC;^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):"));
$write("%s",("f(\\\"\\\"'Ye%4Rra744(f\\\"\\\",2):f(\\\"\\\"{#tiuqn\\\"\\\",2):f(\\\"\\\"})215>5[qa^32^\\\"\\\",2):f(\\\"\\\"})959(f\\\"\\\",2):f(\\\"\\\"{#n\\\"\\\",2):f(\\\"\\\"})420pY4d8,ba8AAbg8[da304zY[O7bda218lK[wL[j4ldamif+6[ga)91361\\\"\\\",2):f(\\\"\\\"}5[,6[j4lbat(6[(6c%a315133A71/129@31916G21661421553/04[04cva%%%%\\\"\\\",2):f(\\\"\\\"}*+1%%%%811 -\\\"\\\",2):f(\\\"\\\"})48\\\"\\\",2):f(\\\"\\\"{3bhaj:+1 j@34[34cbawm4[m4cl4[l4cbaWm4[m4cba\\\"\\\",2):f(\\\"\\\"{m4[m4cva)(esolc.z;)][etyb sa)t=[#>[j4[<6hea3289m4[x5[j4lba,l4[w5[j4hla!\\\"\\\",2):f(\\\"\\\"})46(f\\\"\\\",2):f(\\\"\\\"{#~~v4[%5[j4hea(rt.o4[z5[j4hba)A7dda\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"};l3efa~~dneo3hra~~~~PUEVIGESAELPnr3ala~~1,TUODAERw3a63j$a(etirw;\\\"\\\",2):f(\\\"\\\"};u=:c;))652%%%%)u-c((||13jda#-<q3jda||i)3mhaBUS1,ODs4qka)3/4%%%%i(N4cx5kU4xPa2=:/t;2%%%%t+2*u=:u\\\"\\\",2):f(\\\"\\\"{od7 ot0 yreve;i-=:u;1=:+i\\\""));
$write("%s",("\\\",2):f(\\\"\\\"{od))1(evom(dro=:t elihw?s;)s*45oi5vv3jd7dladohtem dne.s3dganrutern3d~aV);gnirtS/gnal/avajL(nltnirp/rZa|atnirP/oi/avaj lautrivekovniJ3d.4j[2cib\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"};0=q;)]q[c=z(tnirp.tuo.metsyS;)0(tArahc.y+z=]++n[c;y:]q[c?n<q=y\\\"\\\",2):f(\\\"\\\"{)0>2%%%%++i(fi;48%%%%)31-)i>3c&as(+87*q=q\\\"\\\",2):f(\\\"\\\"{);41122<i;(rof;n)rahc(+K4r[2k*3&oa=]n[c);621<n++r4aqa0=q,0=n,0=i tni;N3&ic6ayi4asdRbQeslxfvfllRf<bedRb;f<6;agb-a|dzdxdRfGb8aqeRdYd5aN1Gi;agb-epb>aqeRdHa>aJaRaAdteFbaeIfOa5aEg9Y6f9aVG4aLa7a;a4a<aPhsmkdxd;aNa?c6a|eebHaFaIaebzeJaeb9a/a6a2dQbUe-f2a-f9aVG5d6cRbC3gYc-f/aof0fRf>p5aIh5eZo2e6aRa;dNaxbogj+Gh;aTapc4aLcEeyiof6amc<byg-fJlsbvh3pWfybxcxc>aGaUeAa2a6a\\\"\\\",2):f(\\\"\\\"}g7a6a@a\\\"\\\",2):f(\\\"\\\"{g:a?aMbKaKa6a?e:a@aEa2a|gZ"));
$write("%s",("fMbbgli>a:b1a-gqmUf\\\"\\\",2):f(\\\"\\\"{bHa4atcEiYz1j3bD1Ec3b\\\"\\\",2):f(\\\"\\\"}bJaMa\\\"\\\",2):f(\\\"\\\"}bJa|UEc-bJaJaUa-bJaMdJa8bKr;a8bs-Ka8bs-LBwbgMPaOaNtYz9bKa0+P|Ta0+0+<pYzYCJaLaJa0+;ph4eoa;p1MYz:b+b3b+b(4akagMJaHaJa8b93a-aHaJaFdS5;a0+Ua:aUa:aKrviSfQfRl4al0sbsb2be3^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'maviDa-a|bV2-a@6aua?aGaUe>a5j\\\"\\\",2):f(\\\"\\\"{gKaKa|gZf~6cgaagQjkg&6esasbvh*b-a/bxcHa|fNke3c0c\\\"\\\",2):f(\\\"\\\"}b\\\"\\\",2):f(\\\"\\\"{gph\\\"\\\",2):f(\\\"\\\"{gvg1a-g\\\"\\\",2):f(\\\"\\\"{bHaNkRf-e:a:a\\\"\\\",2):f(\\\"\\\"}bHa?a\\\"\\\",2):f(\\\"\\\"{gJa\\\"\\\",2):f(\\\"\\\"}b5aAdte@a1a-g0iNkxcpb7anb2b:b\\\"\\\",2):f(\\\"\\\"{g2f@j@d-aIfekx"));
$write("%s",("cHalgjghgmk-aUf0ixiRf-f-gSf|fNkzeSgxiHack;a/aDh<b+hWh<apb/aDhWhnb<aoI:b\\\"\\\",2):f(\\\"\\\"{g/aDh-f-g+gFa,i|b1ali3b:b\\\"\\\",2):f(\\\"\\\"{g9hHaNkHaUe-iCe|bxc3b0a:b\\\"\\\",2):f(\\\"\\\"{gIa|bzeJa|c5b#aQbxi<b=a-aHm*c3bxdUe=a-a?arw9ai3eta2bMa7arh|bphnhlhjh9m3hAaAdMUPcgfvfOhJh7aEa|b8k6kMaHm*cEc,dJa>a2aIfzjMgMa?arw<i+cbi6a13k[axdtbg\\\"\\\",2):f(\\\"\\\"{8g/aDh=apiRa6?Cd6?kb-LXa,hDhsk6a7b5ackRfwb\\\"\\\",2):f(\\\"\\\"}jUe2b5a9gYi4b-bhcxsOiOiav0c/bxd;a<hoj-?aea6a2bT>cwchKZH6a5n2a5awnQT\\\"\\\",2):f(\\\"\\\"}gEhgl7tOi6aUhvnHa1dmdLhRfXkJkHa:eXkJk;l<b3bxd6aIhDkPh4ljbkikixb9iacPa;a,bOhn5fbpbubld1bZb,VnbpgujsjiiR3RiWkuhUk4j<b<b<bFj:b<j<b<b,cKjHj7b-bKjEa?aSg3bDd0kMi9a7b6g-a5be6,cKj=a9a7b.Aq3e33gcaCj33eea.b8fE3c33gfaJb7bdU3fmagkEaHs9aH/xbu3amakiykpjCk,cKji3asapmhh.bfh,cKjsbHa\\\"\\\",2):f(\\\"\\\"}g\\\"\\\",2):f(\\\"\\\"}5c^1"));
$write("%s",("^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'aVjDjCaLi6aakflhk4j6aKk8jYjel.k<bzeSCc93gca;k53cEaIkGk3a6a<bkicjPT2b2a2aWRekZk0iwb\\\"\\\",2):f(\\\"\\\"}jRfhDnc:e7b5aWf=aKc<z\\\"\\\",2):f(\\\"\\\"}k5a,bJa6agAa%aub9h5aUgwb\\\"\\\",2):f(\\\"\\\"}jHa:e-b9a9b9apkekyg>am3awa@a@aekyghD:a|b9a0b9ahDNBamb>e|bPg9bJa0bekyg-b9apk9aCaAaJa9beknbJa6a|b5a,bRf:e-b5aintb-ajh9apb\\\"\\\",2):f(\\\"\\\"{iTTDXviWRyg8bAdGh-aWR*bV1-aWRyg7s3h13ahbXb;d9f/bxd6a-b9a8b9a7bJcJayb5muX>aJa*c@dxc?bsuki>aJa-bIlteUehDR2Kd/-vb:atcJaub5aEcxbR3,b4b-bVgg;aiaTkRkmdLh^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9)"));
$write("%s",(":f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'7gycdlblpb;awb\\\"\\\",2):f(\\\"\\\"}j*l3\\\"\\\",2):f(\\\"\\\"{aQ<ZE<TTZHoM;ZJdHd,l2nInClmm9n7n0nG.<nD9hbH6Ar89;uVvMVMvHVIsEa\\\"\\\",2):f(\\\"\\\"}bDaBaEaSxubvvlbr-t\\\"\\\",2):f(\\\"\\\"}6U|bs-a:t0\\\"\\\",2):f(\\\"\\\"}|r<8VUn0*z.09Unfbiws0uvhxttio5bC\\\"\\\",2):f(\\\"\\\"{gb9bZ8U4L6hb=aD9hb?ak:EavN|RHkA9@afb2bib9bAazoCr9DJ|Qp\\\"\\\",2):f(\\\"\\\"{ia5czdGU3HkbU/Io1<Ea5bCy6C*.>ws1db\\\"\\\",2):f(\\\"\\\"}b,oTRWacphb3bMo=pEE/Keql\\\"\\\",2):f(\\\"\\\"}CwU8DrN\\\"\\\",2):f(\\\"\\\"{Q:fw?sn3g5eQdAZrC4Z4Z+5E>t?4p3|w\\\"\\\",2):f(\\\"\\\"{tj,/bN?,oq|Tnjb8baRYzUiYa6XZvCyOq|bXo?/Wa?azYD|4VykVv.b1bq\\\"\\\",2):f(\\\"\\\"{eDkbAo.3qUrg?w?aE@l\\\"\\\",2):f(\\\"\\\"{tmF1wbM|vbW:hxqxo+?87|\\\"\\\",2):f(\\\"\\\"{bS4zt<yjbq+Xa?9rDq|\\\"\\\",2):f(\\\""));
$write("%s",("\\\"{BcKnoXafxA8g,p4I\\\"\\\",2):f(\\\"\\\"}Ezt?0|pGn:8bS4NazWJ\\\"\\\",2):f(\\\"\\\"{-jdb\\\"\\\",2):f(\\\"\\\"}90x69mjNaCajbP\\\"\\\",2):f(\\\"\\\"}6bpq\\\"\\\",2):f(\\\"\\\"}F3HWaCa&6e*dDa6o0rzbKubb-jB39FM4<<jbTp<atK-1XVS\\\"\\\",2):f(\\\"\\\"{Qaebvb9bDaQVSa20hcy|=9,b=BYgCrvY3vZr89QQebY<7blbR+W8n3/bZtTo\\\"\\\",2):f(\\\"\\\"{b|b<a5,M\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{t-b9IDt-dyb5D?atbt\\\"\\\",2):f(\\\"\\\"}9Z3Jx\\\"\\\",2):f(\\\"\\\"}VGz\\\"\\\",2):f(\\\"\\\"{p:TaTy|bM<GoROiq,bmsEaYa.l.bB3ooo+ac=HooSzVnlh3JltvN|Rdb7bjbWKFYYadb7bc4*:kYr3jtvxEal@KuL\\\"\\\",2):f(\\\"\\\"{F81>SaZv.bFqrQSaH6|wd\\\"\\\",2):f(\\\"\\\"}zbQpUaAtlb\\\"\\\",2):f(\\\"\\\"}?hbCUEWhblbtUUnc|JKYq38w<=U6b\\\"\\\",2):f(\\\"\\\"{bzOaTU0z0;=a*dhOTTDXK>1:it9CkhWav028uqSxS,S*2EGaVF\\\"\\\",2):f(\\\"\\\"{:po*b|oR>h+wLH6Y.7|nC|oTax.Ta4qH63b7T424T<o2T4bs-EaEwEqZteqjbFmtRMoDa*xc\\\"\\\",2):f(\\\"\\\"}9blWtRvbuTVa-pFT*.hTkDN"));
$write("%s",("ab.ZtjbCaFTurk8*.t+uqQ|b.\\\"\\\",2):f(\\\"\\\"{be6G5x\\\"\\\",2):f(\\\"\\\"{6rSSkbzOb1ArVDj,o2Z\\\"\\\",2):f(\\\"\\\"{b4?rpo+>G5Z\\\"\\\",2):f(\\\"\\\"{<OSaGrEwjbDvs1fbFTUaX,*b+bG5e6pohb,b+re6G5sqAoe1++4bSajbFa2bD5b7zO0b5bl9OOlbBaEakiXwkbDa7zH2lWhPNaH2b:e@bEaEqq.++|oEqe1++jbvo*oAnKz<-I/1b6X;<MR1bgb|?=r-bPrOv3hmY7F9oOpVaki=RhP:Rgo7R=aTa:6NaCa26Aq0Ry|8.+|i\\\"\\\",2):f(\\\"\\\"}TaJr|RpwZa?aDa*b\\\"\\\",2):f(\\\"\\\"{rDavR7F+b<a.5hb:W+bhbdb*M/puqo3cyaNa7F2MMwW:KrhbP|DaEyzt=a%3eqbD6eWR0TpPQ=aTaj+8obs?aKrhbPv+3:Wqveb?aCp@a4bHk/R/=4oibGoLpP57bR=kb|b|pzdsK=WHYM8lQTYEahQfQfpdpybUa6r*bLR@f&dNajp@H-0Q:9fDa?/MR?aPa@;Xa0bW\\\"\\\",2):f(\\\"\\\"}p?r\\\"\\\",2):f(\\\"\\\"{xyRahbNaxwLBsvW.t>Awz*S4u0I\\\"\\\",2):f(\\\"\\\"}bbjx?sab=aTs+b<ao+Tp4Y<ao+hbx2K*m|vbluM\\\"\\\",2):f(\\\"\\\"{mb;ww;@aDa*rlhnzlz<<1xsz<.>aNY9D?aMROj5Q.7ebA?Y?jb8b\\\"\\\",2):f(\\\"\\"));
$write("%s",("\"{Atb\\\"\\\",2):f(\\\"\\\"}8ebo\\\"\\\",2):f(\\\"\\\"}t\\\"\\\",2):f(\\\"\\\"}gbk-pSXoiPluebo\\\"\\\",2):f(\\\"\\\"}mb8.\\\"\\\",2):f(\\\"\\\"}SiPEa6+ybcb7zJoIG6b/bdbhqN\\\"\\\",2):f(\\\"\\\"{</abJoY?tbXaCawb+6.KP+66vYZa:-?GOa1511Nv<3uJiGTay>CoQQlPybPa?|xZ6fS*Zb./2b707p,\\\"\\\",2):f(\\\"\\\"}.6e|dkbslz5OjS*ubLH<a4b8,@22bX\\\"\\\",2):f(\\\"\\\"}W3uby4DaUswYatYoP?iS.M/beqibVaDa9vH6vREtl0iP-:fbgbJd++Uaebyb0O?6O*@aS*fb98?03hh|J1p1SacWhq\\\"\\\",2):f(\\\"\\\"{O,vjbl-8;Ds67dqB|ATfXtMWoRxS00bsmIwnqQaD-2\\\"\\\",2):f(\\\"\\\"}fbS*twCa|bSz0x+*jtDaS*2B:t1jXi:\\\"\\\",2):f(\\\"\\\"{UaYUk0+bcbWK=>OhFa<>1jYax4Buc,\\\"\\\",2):f(\\\"\\\"{3FaaT\\\"\\\",2):f(\\\"\\\"{*fbo\\\"\\\",2):f(\\\"\\\"}T|P*gbXtVabm2bn-ATfX+bjzzYEjKYd\\\"\\\",2):f(\\\"\\\"},b3G8;6;\\\"\\\",2):f(\\\"\\\"{SYAYa1bYAkiXw(6e*dUa6Wzb6WOa/-tbybzbG3fb|b.dybBa,9t0Hd7bHQtWsoNao+JsM*|bPsP*gjeFyb7VYrSrT\\\"\\\",2):f(\\\"\\\"}eb@>Yai,Asn4WU?0"));
$write("%s",("|>?vuynrQa-bcbfbNaN1c\\\"\\\",2):f(\\\"\\\"}v=|TCGSa6qv|<UebI\\\"\\\",2):f(\\\"\\\"{VoKEzuQP*bO5V|kbbD+U0bWDn-6rN0VF9bnoKtI=zbnHtbTEa-mW0b0O\\\"\\\",2):f(\\\"\\\"{bLUbDGFV?\\\"\\\",2):f(\\\"\\\"{b+2Faxqv3pXByXO9bhb4udb9bQqOqcb8rl\\\"\\\",2):f(\\\"\\\"{RJGM+U0bGpzb?aebybj*8;|vdb;idpoSuLBZN2wY3b\\\"\\\",2):f(\\\"\\\"}btb20Zl23yb=a0\\\"\\\",2):f(\\\"\\\"}Yars6WE0Xs(DgpbJViPAn=|zbVabm5bawMV/Rv5W.Pa9,7,Qr3*yb<aQ,.bVa>v8*Ts27M*K*YaXsebS*ZaZalt\\\\\\\"\\\"),\\\\n(\\\\\\\"\\\"1bvb>aYzlTS,s<6zL\\\"\\\",2):f(\\\"\\\"{kHZB5QG@PaxZ^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'3elco\\\"\\\",2):f(\\\"\\\"}d4f\\\"\\\",2):f(\\\"\\\"}VaS*.b@,zbv\\\"\\\",2):f(\\\"\\\"{Aa*\\\"\\\",2):f(\\\"\\\"}tK+y|beb9b<1"));
$write("%s",("3Tw*ibAIG5PqefAa;P=Bq*o*6Y59YMxhczhp857*:,..Oz6blycbEa0xW\\\"\\\",2):f(\\\"\\\"{pU1>csR82W2u:tjtht|bNaTuYp3bybBaO46\\\"\\\",2):f(\\\"\\\"{Uao|1MeI\\\"\\\",2):f(\\\"\\\"}Q381bjb5bGp0bkiL<zObbp4p06-J1tb3trU7bxrtbLp\\\"\\\",2):f(\\\"\\\"{LEMU1Kf$dMhrzDiG+Mhrz*t1bu,>00Fl\\\"\\\",2):f(\\\"\\\"{|QAa7q?sybPaOz1bdzp\\\"\\\",2):f(\\\"\\\"}9bNaDv/tabjbk,bO8@Kfdb@2ebf-mbNEgb,\\\"\\\",2):f(\\\"\\\"}.s\\\"\\\",2):f(\\\"\\\"}z*ti1|Ud,a.ybcbKWRLldb2xtZ|kbmb\\\"\\\",2):f(\\\"\\\"},X\\\"\\\",2):f(\\\"\\\"{boZtybzJvySqBvn:hpq:Bvki:y.bL\\\"\\\",2):f(\\\"\\\"{E@KrdKCw80@aki*CD5Qakb92vb72qrJ*UrX\\\"\\\",2):f(\\\"\\\"{k:aq,?3bz4r>v-|bPyczjbsu2EkiDP?sybj+vC@qykybwbibzIm5M+LOK2=|xOCCR82ug,-pxbhb?an:,W\\\"\\\",2):f(\\\"\\\"{Ac\\\"\\\",2):f(\\\"\\\"{37=Hz?<a:\\\"\\\",2):f(\\\"\\\"}rNvV5bW,fbuu,6e3ay47kNa?1kbv*wkSq1,:xBaO|z:?aO8+9Va12mbOO:,:8JOb8clbCa9u=.Ta:3cb83T3H4-LF\\\"\\\",2):f(\\\"\\\"{/4H4Ua?s=*Znp0t"));
$write("%s",("b*v,*2K1b*bR8kb1F9rwM1:Sz0xUza-SyEa<tfG1zXargvoJpmVgbIr+LWX5bv>a2bbDrwW1x?CaOJgNixtb=aScKZhjiw/\\\"\\\",2):f(\\\"\\\"}/*>aYzhbi-N?fc9bmjHqPa7|42fwtbNyAoVq?pOG9Gz?tbtbog0b4bVaMCai1:yb2zZE7z@:gEU+8b<abbeD1:LSfbwb>ipy/bs5Xq*6eVbubx\\\"\\\",2):f(\\\"\\\"}R3C\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"{*DaU1r:jbUao+Aiab9Ki:=xi:S79f4bub\\\"\\\",2):f(\\\"\\\"{*DaLG<94bBvjmn7P5?0*:Aav*Ut\\\"\\\",2):f(\\\"\\\"{7y7pXS0JzjtUr|fVa37qNQsbboZebub9ffb|b0.WabqX|urF.|VpEfpI-\\\"\\\",2):f(\\\"\\\"{rjb\\\"\\\",2):f(\\\"\\\"{beq2br.Q,<-N|VaO|Q7-pYSg?F....OwbcbX>a$bvbXQv*<38rhpiTP\\\"\\\",2):f(\\\"\\\"{r8t0?o5Mt,XoVM@/BuBa\\\"\\\",2):f(\\\"\\\"{<-8P?iD|zB.VaWa<yZ+Z-bb4ElbSazbNv6qv|YGasZauG**F5GMwYY9W9gbXae?N2wYZaEa5bXaEq-6WD,6exbzb8babtzV5Eagb4vtb4b\\\"\\\",2):f(\\\"\\\"{=zt4b6rlW\\\"\\\",2):f(\\\"\\\"}KAakOHJpZ.*4t:\\\"\\\",2):f(\\\"\\\"}Xaarj*4BApV,AxUr?Cb\\\"\\\",2):f(\\\"\\\"{9*Dz"));
$write("%s",("ub3;ki1;fbu|tbAakbbtSaR=Ya<aj\\\"\\\",2):f(\\\"\\\"}Pq</g5\\\"\\\",2):f(\\\"\\\"}EJ/<:aacfty*+b1:+XsuO8.p5?3buynr7Q0t=Bibit\\\"\\\",2):f(\\\"\\\"}b3hmYzq5?\\\"\\\",2):f(\\\"\\\"{=87rXMlVwT:g5\\\"\\\",2):f(\\\"\\\"{bXQRL2xdbMv\\\"\\\",2):f(\\\"\\\"{=SxW8fxj0,?yxz;LUMv2uEsq<Jy<aRY/RubQaFazbq0PXQaDaOvR6h-3xl:AoB8g?B8g?OzoB2blT80g?Rn-pUzbo9+0botlb|:Uzz4#Kgzd0W5*lD\\\"\\\",2):f(\\\"\\\"}-7vkbMs.A<LRaIqyudXs.|beb7|9xlbfb,CUa2gD-\\\"\\\",2):f(\\\"\\\"}k2hkbiD0.CK>*=aF\\\"\\\",2):f(\\\"\\\"};O.FwYj4|wk4OGCCOEKDY+g?*Yr-@yF\\\"\\\",2):f(\\\"\\\"};OR>kz:vnv<LWX4-8tR>OaRRb\\\"\\\",2):f(\\\"\\\"{Gqki:ym=X67bL\\\"\\\",2):f(\\\"\\\"{wCd,xos/2E7C|bfDFa2bvbIAryo?56R>.0=HNaG.NaEaJ.+Ehb7F-.Xas-Wabq=aApbb7b,b9bcbUBCxxr5Vw;\\\"\\\",2):f(\\\"\\\"{t@aAIHEPqOz6bJ8WYc\\\"\\\",2):f(\\\"\\\"{AoiywwRx3x4skiGZ;,j9<*9|@i|b?GvTuLYg=u<a,bKGe=aZHoMf65z.=P;-p\\\"\\\",2):f(\\\"\\\"}90wGyS*ubDtxbQ|Dr|E:t\\\"\\\""));
$write("%s",(",2):f(\\\"\\\"{b>q1hfGLwGCcbAobTAo%3c@bNu?QJ/ab/R..e?Pc\\\"\\\",2):f(\\\"\\\"}>vvhbOao.\\\"\\\",2):f(\\\"\\\"}r8*tB7=FqYU?v,b8b9oVC6;Yahv;q<L-bDsgvo.lb>a8*\\\"\\\",2):f(\\\"\\\"{bR8?*sB@vdzZqk+Fpr-v>Oao.hbEq@vU>3bb\\\"\\\",2):f(\\\"\\\"{g2S>ub7;o+HJ7o\\\"\\\",2):f(\\\"\\\"{x?a:sOA*+e?y92v4B<w67o3cQaPvFa37=HWDj35bPv7=zbKGmXOrnxC*nxB3iDubrQS+k2?+dbS,EaUa=aeyo.DaYaks7b7gD\\\"\\\",2):f(\\\"\\\"}GM-FS9e$bBazt,bBN/b+bfWG@X>9xb1wYarJBKsc\\\"\\\",2):f(\\\"\\\"{y-uyVP6B.bOrkxbV.b2NWXFuBq?a*+jbFu@a>qXt9*6qZ+Oa7bhb1b,jLR\\\"\\\",2):f(\\\"\\\"{+@xfymb/y7bvXKsZFYa<DQQjb6;i3cSb+bboxY-.?*bV6b/ykxjx.Oabebcb|zPaoyGMiqUB-bKTfbcbgvebvbfB<sVVKM2z5bhbTuvfOrQsS9VY.bUpTu2bBG6WzbdSy-2ztb<\\\"\\\",2):f(\\\"\\\"{SqzbKvX\\\"\\\",2):f(\\\"\\\"{H0ZagWn:|vdb7brsYaybP\\\"\\\",2):f(\\\"\\\"{s\\\"\\\",2):f(\\\"\\\"{|vdbqr|b=HBfzv\\\"\\\",2):f(\\\"\\\"{bwvM@ku\\\"\\\",2):f(\\\"\\\"}v:JccA,6fac|=arIg9?\\"));
$write("%s",("\"\\\",2):f(\\\"\\\"{bCaF|ure-u,*b0b2zDSCGacpZ|,wvvf3r3b@hZQr<.w<sBaO,AIe-=aXsJB6Cr1Jqjb@\\\"\\\",2):f(\\\"\\\"}<aZ2ld1bb\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"{bIq8uZaCo3b0L:/+ENabTp+nG1pq:LyXO6OUadG+r\\\"\\\",2):f(\\\"\\\"}rAI1bYA7bLyybgf@ayb9sNK>tG?bkv58xn:PrFa\\\"\\\",2):f(\\\"\\\"}b4*i3atbTE@.wb@adkNabx\\\"\\\",2):f(\\\"\\\"}b;v\\\"\\\",2):f(\\\"\\\"{dUad3?aQc+S-bxv6zlu:=Aaxjo;du8bG?btfhYo0+9rYaT\\\"\\\",2):f(\\\"\\\"{=aAnp3cbfb/KWLxvUaO;efhbSag8<9abCC\\\"\\\",2):f(\\\"\\\"{umbm|&6ezd-r,bv3n;y;pyBEcq>avyAostx9hb3b?aybcbOjcbZ0X+\\\"\\\",2):f(\\\"\\\"}kno4bvyXilu2=b/ru\\\"\\\",2):f(\\\"\\\"{th-d,h-aTykT\\\"\\\",2):f(\\\"\\\"}I\\\"\\\",2):f(\\\"\\\"}Z+*=>a,/GaqXI\\\"\\\",2):f(\\\"\\\"}+=ub\\\"\\\",2):f(\\\"\\\"}=\\\"\\\",2):f(\\\"\\\"{=k\\\"\\\",2):f(\\\"\\\"};@3bxtWaZ-/.Oa8pCq7|Paj+6TYgT\\\"\\\",2):f(\\\"\\\"}LyX\\\"\\\",2):f(\\\"\\\"}gqp3\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}Gac=Y-p;u\\\"\\\",2):f(\\\"\\\"}qsOavy9<y>"));
$write("%s",("4y:-.RiyabRL3GFU/R1b,G?wQaz:<;jbfz6,Xi9bhb,bU8\\\"\\\",2):f(\\\"\\\"}b>ihTub9-f8wByd7bmbz6>xQN*bGo=HdWgp0zub9-lvmOb/p;QqQaFa1:?4W857-89bhb5bQa571b&6e/adz/scJ/=Wz<0jw7bZa\\\"\\\",2):f(\\\"\\\"{3E/U/eoM7hbdb=BBGq23IC-1Eeua+GVKRa|bE/-|SaQ^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^32^[2fha\\\"\\\",2):f(\\\"\\\"})3(f\\\"\\\",2):f(\\\"\\\"{#v3mja13(f\\\"\\\",2):f(\\\"\\\"{#,4353(|a3891(f\\\"\\\",2):f(\\\"\\\"{#(ntnirpn\\\"\\\",2):f(\\\"\\\"})4201(f\\\"\\\",2):f(\\\"\\\"{#)~4[~4bGb7Q?Wy?a:9izVavI2b.bBZh+l;xbGatXO5z21hwbjJQ-\\\"\\\",2):f(\\\"\\\"{f2Embvqf@v@BZfgFxlP+Fq@4=KvbbF@9@Ra=Iz\\\"\\\",2):f(\\\"\\\"{izVa7@f-CvL;l0wW0+AQWa7bI-JKY\\\"\\\",2):f(\\\"\\\"{gbbbTavjinE\\\"\\\",2):f(\\\"\\\"}iDKATaZ,U2v@x*BOE@FJq;xbYaUaI3aEabbZ-L9Va3brs8tdbo??fNaS5xbAoB@wbl,FJq;2@v<E\\\"\\\",2):f(\\\"\\\"}5|866bkFv=32|bs@UaQ-2[g^1^\\\"\\\",4)"));
$write("%s",(":f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'d/dGatXu6RaWa8Imb<=D*\\\"\\\",2):f(\\\"\\\"}b7@3wWa6H-:GtjA.be?xtz-Ba|pA|?03hh|J1o?Nv2hCpQazb=.z=Pa62|b=@LXdz1FTac.<Qcba7/Kk43\\\"\\\",2):f(\\\"\\\"}-b@aQ,+bNargaPz\\\"\\\",2):f(\\\"\\\"{WwPNz9SBuyPa7SOtG9dzBY=|7.rgTEFvH/,b6qDaEa<rDaEPfbwbz49Cjb2bA+Y>1bh-z1jd:@<=a<y-S+BEkiGZA|zb8uZaEi22=y\\\"\\\",2):f(\\\"\\\"{bl85QK5mbg|*bqoWK4IRq2b44ntcbabv@ai9H+W6,./du?a9t2bur*w8qi7P6kWpjRaWadAX0[f$bmbq.q,yuAaj=Vaf.S*VaWagv@aP<s-Wa.bVa;<l9RarXL<VuUa5v/K\\\"\\\",2):f(\\\"\\\"}QbmFp/ydKCwE:EE3v.OfU|To2BaCab9./WaW9n+6b@a7Ijby*yCTsC-aboZiuzbz4c&b>Ijber|EUt.b>qG@Ta9rdpTaBqywkb62jy*zQ?Xa1Ho|xT9K\\\"\\\",2):f"));
$write("%s",("(\\\"\\\"{b|biq6;XttL8qUMyb9*fb12hh+bhb1x=Cu=*zWKSc>0.tbboZU3QadU3b9QVskbvXQa3b/DF4e-a27Pa<3rQ,4W-cb3gUDcblyp36g=@865Em.<2b8Or06e?aaFLUVaebtoVa3:ZO90|yDasRe;F*y7uye?zbapAq+bXVSQ\\\"\\\",2):f(\\\"\\\"{bh-koUY/YG/JUcSal.\\\"\\\",2):f(\\\"\\\"{0lbdbx+HoGaNW\\\"\\\",2):f(\\\"\\\"{bjbO8j*U?Kq=HOzq1q\\\"\\\",2):f(\\\"\\\"{SQ|vDxLyQa+bgv1zS8CFDa,w8.abB;W.*+K7ufeqoBK3csa2y:9/|@hX|DF+bAaN||Ua\\\"\\\",2):f(\\\"\\\"}b4Bl+zSB;zbKGk|Y\\\"\\\",2):f(\\\"\\\"{tRKMxby>cbcbr<7=FFH4gw5bzb6b/biD+G<J=C4;?Xjb\\\"\\\",2):f(\\\"\\\"}>cbEaKvU4ZaYaHpaxDU:AZaPvur2gu,mWGaVFg4TadbcbgvTR\\\"\\\",2):f(\\\"\\\"}Fd9j,Cfqamthb-bQs@a5x1,Fu9LaM3eyapXSaTR:Ahb:s7Fko3ZDUIgzvRIa.b?92bqIFITa,IGam8Faj>h>,te>iwqrrK,b5=Pq/tnB|bEaYa>s.wCq/b/bm+Ya|t>a9IQrAw72=awWVamb++F*Saqzi/Dz40.q<ad0VaAa.-+d9?6UE0?|yx53kbCrH4eHejbvj@a@aDp<L,,hb\\\"\\\",2):f(\\\"\\\"{bpslb?a39Bq39ibcbD9<Q1"));
$write("%s",("14=lb.wd+3x44ybDH9g9bH6zYEjKY2>=RjC6FbT;<U+Yrz\\\"\\\",2):f(\\\"\\\"{vb37Va2JBaWy06ezdr=Tp9b|pb<n4eIFI;Hww/-dt|Vub1bhx@aE+B\\\"\\\",2):f(\\\"\\\"}i:\\\"\\\",2):f(\\\"\\\"{uGMjbF+Wa>Eix9b<aQ3Na@hEaiG4bQzxblbmo2Ouqvbt053lb;qufmo.OQzAohbH6rKwb<r4,F5dW*oqHB;KuYzA6@2Sai>Scu1DawMo|/z/6/zHwDwS+3b7vRnl.|bgvmKgv58mb>W|b1FSa48xK<9Va58Dw5=q-D60.aFubQa3bab0.,bo2e-ab0h<90hhwSrnG7vX2xK\\\"\\\",2):f(\\\"\\\"}<Ya@2DwS+AIB+gvlSQQmW4LKsT-z*k2v5Dw5=7tV,&6e?a85@2Sa5pHJ0rtY6<q+XaU885cJbb;T|:xt|:,3F\\\"\\\",2):f(\\\"\\\"}mOTo6b5bH4P2|b4bwwe3qEa|>|oR|Pa9gybPa9g9uLpmuQ?7;0bR7lD*bdpRL7SmoM+Z25,c1YhyMfh+zGz4\\\"\\\",2):f(\\\"\\\"}8bB6a=bbbUz11OPYadk;wVuB|vrKvw4Faab5b6YF5ibYaF5a\\\"\\\",2):f(\\\"\\\"}F5ib0bDzDwJCv|cJ9fA1c2bb-qw\\\"\\\",2):f(\\\"\\\"{koCwAoU:u.d\\\"\\\",2):f(\\\"\\\"}IUu1dY,bMzzwF5B1fb4wxb*o65*b8qw\\\"\\\",2):f(\\\"\\\"{;Kjb9K5bNuK*:utbKwty=/yb"));
$write("%s",("<K2b/^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'=fzdS5;s0Ds*xTYp2x2hm,Yp\\\"\\\",2):f(\\\"\\\"{bLUWXYaIdKW0b?4Qx<aS+|UKWi9zwut1AGQ?vcbL->0\\\"\\\",2):f(\\\"\\\"}Qo,YSBaW16,/sFaQp6b9*otDp<=l\\\"\\\",2):f(\\\"\\\"{,bX55Qv3pXH6NapX9b?aW36,QazbX=1,Qpogc\\\"\\\",2):f(\\\"\\\"}o;dbXt8:Zn?=D1F*gbJ1Ba*Iwbur.OOaO8mb9L6X*+z1L;O*btS2|J;9GgabOj>a|Ul\\\"\\\",2):f(\\\"\\\"{U>aH+bMLIdaJ7v+bCptw<aVa;rfzhMgbn:hbYAFv3bU>aH;rYN-bUB\\\"\\\",2):f(\\\"\\\"{u0b5biY*zabAy<K6?jb4-,b<a.=fbjd&6ezdfb>at,Fa\\\"\\\",2):f(\\\"\\\"}bj*ebzMMw2xcJ4rauXy*+z1/C59/DVaCCR8b2Wy4-OG\\\"\\\",2):f(\\\"\\\"{On=ybRa<,eF28mbZa9.o?/RzbU2B16,,bM0\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}PacbJ.L\\\"\\\""));
$write("%s",(",2):f(\\\"\\\"{70fbuGmb-8:I<*\\\"\\\",2):f(\\\"\\\"}b|bZawYyHbY9qab\\\"\\\",2):f(\\\"\\\"{b4vtbvqMLAaOHMHTD|b;zIz<\\\"\\\",2):f(\\\"\\\"{:\\\"\\\",2):f(\\\"\\\"{6b/*suW\\\"\\\",2):f(\\\"\\\"{3qSFnHZaM\\\"\\\",2):f(\\\"\\\"{QazbepQag1q=*bn78b<aVax@:u8QGidzId.rnrc0|oW3?tQaETEaJCjp\\\"\\\",2):f(\\\"\\\"}k1vVvHqt,pEXszHr\\\"\\\",2):f(\\\"\\\"{l@nz\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}Pas2Far:b4jbWar3dzHt8LX\\\"\\\",2):f(\\\"\\\"}oFHy7IoD&6g~bgb4sYadboN3r1Mubtb:Whz2jIQ,jyz\\\"\\\",2):f(\\\"\\\"{BXaNaS,1borb4@a8bQon+LRRKizebSa?=tbp\\\"\\\",2):f(\\\"\\\"}Ua@vWoZQKTfbpNubebSain5sNaAoki:y8|6zb4@a87:vS,1bA3cY22b7F1ZWoEaDaZa7bWaCCkbOJ>|7K2F2+V6KCi9p.|uiztbq.o.9KdXo\\\"\\\",2):f(\\\"\\\"}i>ubiztbybv34xdkiz:uvC2vJRz6:Pp38QnqU89q?07slb:IPVhbSa6rFYaTh2kxa7x|u1377va17v<B7viuKGP5/C2*xZ4bd+i\\\"\\\",2):f(\\\"\\\"{l+8ZTan+joi\\\"\\\",2):f(\\\"\\\"{3\\\"\\\",2):f(\\\"\\\"{QBlMCXxhub+ymovS6WpkkimH2gefJOQz"));
$write("%s",("z\\\"\\\",2):f(\\\"\\\"{6blbCwegTukdNEL=Aoc\\\"\\\",2):f(\\\"\\\"{S*fw0r|lN?S0bbvbA*Cqp7Sz7|qx-b0S7uWY8FjmSY@qPYIt>awbFYFajQNEQagWd0wHEao-X1abw*b5fbS,Ca-Hg|Y0Raz\\\"\\\",2):f(\\\"\\\"{z?ujC-N|5bgviyp40-yPXa9fYzz@?aPVYrmbr<kic+6b|bsKSpVCOaCv\\\"\\\",2):f(\\\"\\\"{bWaub9vRa5x8+CaubiU.7Xy1b4x0tzbabGJu|1rvbTE=a7=vbkW\\\"\\\",2):f(\\\"\\\"}bhb|>I<msKzf\\\"\\\",2):f(\\\"\\\"}Cy9bdbg8hpxy-by-:Jww|9=lqMZPKVCy6bu+zb*<Dig557Cab4?Cu.PaNEI?k>Oa1ru.wLEjvuc|8beqUpyN572+GiFJDi>akiC5|vkiZ7*bd<Ns+b\\\"\\\",2):f(\\\"\\\"{OFIFa6K?hY.?T<y/bzIKv3+wvmogbst.bt:S0gMS>W\\\"\\\",2):f(\\\"\\\"{9Gkip<qj9pwbxq7K5.l\\\"\\\",2):f(\\\"\\\"{>BvU>a2b:G\\\"\\\",2):f(\\\"\\\"{b4r5VRay>wH*,3byNh\\\"\\\",2):f(\\\"\\\"{bbzbjwhwv@bT?q7,*No+RUTsZaLyD9<;g2buywzHAo4V,PLBV6D*kiPUu3W3=a-bXaXi./Do0b1A=aub<a|b2jiG7zabnvlvZ4H6WieImb-b.:\\\"\\\",2):f(\\\"\\\"{xXaWRPTab\\\"\\\",2):f(\\\"\\\"{wTx4BDV/D.s2um"));
$write("%s",("bB/*5?apxS>XSH6jwgHjbAa>tab.btKSadutbiU+ol0,blrWaJ\\\"\\\",2):f(\\\"\\\"}FacqX5GUUB3*Ca6bQs,SzKwH>wHU;42v7vhvOOBv8n<a3O;FVv-j=,1pGam0R,N1o;F58.DzlbLUdbBU7k/bAoOjB3X5DatbQa0Q,bbbb/I\\\"\\\",2):f(\\\"\\\"}nH>a|y,bwbg5rQQS+bkbEaKDGycSh,Gau?nsv\\\"\\\",2):f(\\\"\\\"{ToUr8b;EPawbFJ+E5bbbQyhNB5rQ?tdbR=GaX/z<286,lhcb|bC-@v*bj\\\"\\\",2):f(\\\"\\\"}abB-P;\\\"\\\",2):f(\\\"\\\"{PebGMiGyuQt@lo6pM:liKWRY>ltS*<,>a\\\"\\\",2):f(\\\"\\\"{SuqpJ+z2bbbi,q19Tybr<-95|5E|zxtq;\\\"\\\",2):f(\\\"\\\"}bBpjp@a<1ubT3;s;O+,1jf5tt0S7Kz1vTkbU2nSlSkb2h5gtrlT,S2+j*G/1,.=1|g\\\"\\\",2):f(\\\"\\\"}M+t.|bYomS@a3bb7V*Fa-bcKlb*r-p\\\"\\\",2):f(\\\"\\\"}SE9sLlt5DRa8rmhru-0>a*z3b4rPnQa5D<aQa;O/4tSQo/*5,=t;@M+YAUn+bZa2OW3kipLZ|mLlb<JTa8L|bkb/sxbg?wkUat-o\\\"\\\",2):f(\\\"\\\"}<rFqb7AaHrbS7z2bBpNafb=ac\\\"\\\",2):f(\\\"\\\"{7kmb+9Pn450bXaoobbGF+bWRIbXPhbKR|bD1YaI?NHa9\\\"\\\",2):f(\\\""));
$write("%s",("\\\"{<9DubYaBE=rm<eq69vyYo|8Xyhx<J2:D5bbgbq2hNv=1b-GItY24btl2,4vYMubzt,o:|ItJrAaYa6z0xhPpwP+QahxjbybAJp*AJVM3@7HX2YNWQ?\\\"\\\",2):f(\\\"\\\"}Hy4LX:izbcin\\\"\\\",2):f(\\\"\\\"}ztb.bk81bEQZ|pyIt+bl2Xa@AItPav@Ga|74wPa6o2b+qCaJqOa+yUa\\\"\\\",2):f(\\\"\\\"}9Farwl0ebgbdbwJQalbKDgb+beD@a<pS*r,B.u7R>4\\\"\\\",2):f(\\\"\\\"}?0Za-b;tiI*ATams=vXotwCwlb/br3<pvbnq4qjm9b3qruXaCF\\\"\\\",2):f(\\\"\\\"{b\\\"\\\",2):f(\\\"\\\"}bXaavS@PBL3iO4bS00vVrTEDIdbkrm,XOQq53AyQz0FX\\\"\\\",2):f(\\\"\\\"}8OfbAoFa5qt?s-jqfxYqx+db4bzbyP8bJd6?B;Z2nrGpd<OGAp=G;2GtsFRoGMOzg-e-a<bb70ubr4M0s<m?bbOwubW>p3wb0yd,gb*bd,;>egLo9d=aeb,br|6bIt.jj\\\"\\\",2):f(\\\"\\\"}-bd\\\"\\\",2):f(\\\"\\\"}gbl<Gahrs=5oz6j=:t.oD/372j7F9b>a|b-tf/4u=>\\\"\\\",2):f(\\\"\\\"}24bAaNEWzhNG2?ajoF3\\\"\\\",2):f(\\\"\\\"{O0bS>hb2bDadbB\\\"\\\",2):f(\\\"\\\"{o\\\"\\\",2):f(\\\"\\\"{Ry<F6+Sa>a67VaZp.w8n6rPa3qCp5+3+xjXaxbNa8"));
$write("%s",("lgOspgKYCawcAeDlbU\\\"\\\",2):f(\\\"\\\"}Op4bt|f>t.*wN99-I:dbPa\\\"\\\",2):f(\\\"\\\"{L\\\"\\\",2):f(\\\"\\\"{bCx\\\"\\\",2):f(\\\"\\\"}Eht/z57dbL;0NJ?S|rN9b+qj4zA4py?y*c72,d|:A98b9-Gyk-9tb=@n9d5cw@z<L/-ZanGQ?Nw>agb87Lo+bQofb87?a1b5b\\\"\\\",2):f(\\\"\\\"{bHtn?gbvx@\\\"\\\",2):f(\\\"\\\"}Cxdb3bFH3gq98-Oas,A*0b?*<yUa1b:>9vUap0\\\"\\\",2):f(\\\"\\\"{wp3+y2:jb/bf,-bpxAoP9W587z,+8xKo?f+s<J;U\\\"\\\",2):f(\\\"\\\"}Urk-RLCD0Fvb/bq1f\\\"\\\",2):f(\\\"\\\"}+b4b*bXapy*b>A-6abOGHmK5r\\\"\\\",2):f(\\\"\\\"{Pa\\\"\\\",2):f(\\\"\\\"}EBajxwLRay-i6aIh6C<P@O>PDa*\\\"\\\",2):f(\\\"\\\"}|Zy5s\\\"\\\",2):f(\\\"\\\"}b?0LkRaVG@a,K6HB*8vL05Abs9b0xubk|Wa\\\"\\\",2):f(\\\"\\\"}?GJ-bbk:@?qV<+bs.Ym1<Xar\\\"\\\",2):f(\\\"\\\"{:pP8<<7bl.AwUa3b4;;\\\"\\\",2):f(\\\"\\\"}Sa\\\"\\\",2):f(\\\"\\\"{bZaCt0bMvX1db<au=OAgbh|XaV6S+Hrybw;LJb9Ea<a.bBqNaJKsB6bhDfgJ|?y,.;zQa\\\"\\\",2):f(\\\"\\\"{tUa>qVa082.ib<-67ubDK1b9bl.Vo=\\\"\\\",2):f(\\"));
$write("%s",("\"\\\"{mbW9.\\\"\\\",2):f(\\\"\\\"}v1*bH1w\\\"\\\",2):f(\\\"\\\"{+yjb@A?=r8AIGaqABafbkqxucbQnw\\\"\\\",2):f(\\\"\\\"{ib1bj03b<1>a7bnoZxxbkbrKtbmbvbyovbLsO?ibf-C|+bUafbR=P=q\\\"\\\",2):f(\\\"\\\"{Zavb@ayEb|c919Cai6ND1\\\"\\\",2):f(\\\"\\\"{XH@lVHNG:INaybbb5E\\\\\\\"\\\"),\\\\n(\\\\\\\"\\\"s3Aay\\\"\\\",2):f(\\\"\\\"}H@Yp>ahbc4CtRp1/,bO\\\"\\\",2):f(\\\"\\\"}ix@a-|*bjJzbTaRae\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{b:,zbgbDrRaJ8|w2bR4NalbY4tHN|To4b\\\"\\\",2):f(\\\"\\\"}bcA=H3I@Hi7ybNy67|=Loj*qz=aB1/G*b11?asHwwfbardb=/Qs?aYzUI7b.r:,t0C|n\\\"\\\",2):f(\\\"\\\"}l|DaVaQa@a?I86dz9,rqPao\\\"\\\",2):f(\\\"\\\"}otYq6bcb@HsI\\\"\\\",2):f(\\\"\\\"}j>a=aVa.b3s\\\"\\\",2):f(\\\"\\\"}bWa<aE1SaYa1wP<7b.b1vAa\\\"\\\",2):f(\\\"\\\"{bAaSa7bMq.z3bqIuHGz57Z>iylqxbi?<at<i-0bWaBaOAeySa+y/sAoIrkb<a7bepAa<aIql0\\\"\\\",2):f(\\\"\\\"{b1bdt.bFae;H6L,91R@J,MF=lKFh.Bac|K\\\"\\\",2):f(\\\"\\\"{1y|b72SaOj5bKDCcstqic9RauHAo-i3h=a*"));
$write("%s",("bOaW8cbk.zb@iOal8VaXaYzipjbbt+bibvbd7<a;vrHqH0vMwZtubyb+6S>wb<a5bFa8,>aRaZ8AoDa:s<acbx47zQa9p/lBa7q3zVaYa*b|b*G<aX*IqHm?|dxc03ba4K66bPa+23\\\"\\\",2):f(\\\"\\\"}jmz\\\"\\\",2):f(\\\"\\\"{@q6@1DOaibUau:zbB-Ea/\\\"\\\",2):f(\\\"\\\"}kyCaTa6bS>j97q.l>a\\\"\\\",2):f(\\\"\\\"}GZ\\\"\\\",2):f(\\\"\\\"{c7xbHv*b1bAazbybj,0p<aM*9oAavbvbDpO,E/8rhb.=wb..q:hbP*Ta+7y-Uaty>issuy/lbbl+<akiP/?q2+6bhwL,u8D<@ll6i6NBvv<w9/Za=|iDTu,b.3EC|=/rg|SCxb4bJ\\\"\\\",2):f(\\\"\\\"{lbCaDa+27C*dTClbubkbk2\\\"\\\",2):f(\\\"\\\"}bmbC|ykiqS4=u0*r|W91==aybTaRCDaRaHvW\\\"\\\",2):f(\\\"\\\"}HEv.ebtDTag\\\"\\\",2):f(\\\"\\\"}q9GDU@Lw1bG5q:\\\"\\\",2):f(\\\"\\\"{3wb3bn-H8I+M+Ur.b\\\"\\\",2):f(\\\"\\\"{t7g+oQ,wbgbQygbZatBYpubQoDpFaQ?Y.tbhbibx*yb8.R4|by7+|in<@<;Ta7bjdVaxwP6Y2w6dEj9/bL-,b.bbthD.bc;JyXa+4k0+6h-GtabOCSa5+,b;</C8b,bcbw9>C<C15a-7+\\\"\\\",2):f(\\\"\\\"{dYnIq|bvbwbVaJt3\\\"\\\",2):f"));
$write("%s",("(\\\"\\\"{x8MDOBv/Q@B,ZaPy/|=ro9Pqvb*qCa0|Pa:rqoU3:2ebbbs@hbgb5pa6\\\"\\\",2):f(\\\"\\\"{b\\\"\\\",2):f(\\\"\\\"{*P|dobb.3Za1jbD+8Xa9CMsQ3,/J<>\\\"\\\",2):f(\\\"\\\"{<\\\"\\\",2):f(\\\"\\\"{Lpv.Bufb\\\"\\\",2):f(\\\"\\\"}+/bU:S:9-xbbkNambjw@a>a=s0b2b>w.=Aod9Rz\\\"\\\",2):f(\\\"\\\"}b5|cbmbx*fbUagqGtC-s,wbZ@PmibPaq;b\\\"\\\",2):f(\\\"\\\"{fbBo+xXofb3p4>4bTa69Aa5pmuYp|bg|fbhbz>-jl@*b@aN?PaGrb8qvAo/bl9|v|q:,6b7xVaybOz1p:,X;acr:ry3bYzh,=oDadz9b;t<r..Myl9<rx\\\"\\\",2):f(\\\"\\\"{:qZb:8.b>B+bxhr8avy/N><:O@8bTa=Ah-stL-TzdlU/T3Nkb+Np9bYrkb7bDa.xOaP*fh1v/bWAcbh-Da-qmbo-\\\"\\\",2):f(\\\"\\\"}<VnRaN\\\"\\\",2):f(\\\"\\\"{Jwj2mv?a\\\"\\\",2):f(\\\"\\\"}0ubutabYrH/TaAovvWaN2mbRy>9+odtP*:i|d0Y2lUaw?FqNw\\\"\\\",2):f(\\\"\\\"{1Jr6;bbUyz\\\"\\\",2):f(\\\"\\\"{fh5x=,Ui8gdz1|UaUpQ:F*DaCaVaI<Ht\\\"\\\",2):f(\\\"\\\"}vC*l?9z5s6r\\\"\\\",2):f(\\\"\\\"{b\\\"\\\",2):f(\\\"\\\"}8kb.b1,Q\\\"\\\",2):f(\\\"\\\"{mbKv1"));
$write("%s",("\\\"\\\",2):f(\\\"\\\"}80o;0bpy\\\"\\\",2):f(\\\"\\\"{by\\\"\\\",2):f(\\\"\\\"}ib<wM8xb|bXazb0b\\\"\\\",2):f(\\\"\\\"{=h|4b?ar4B.ab+8ab-7U8ir8wk,6.S+O5\\\"\\\",2):f(\\\"\\\"}bQo2be6:0xrz5WaSa1bS5Qzy,/bmzn?PwNwvni6D,g6v8L>5bSaDaOr-7DyNaTa;@mb5bp;1h7gt00b87WawbfbOazy?aWaFaSaFu4bp;t.wqa@4wi,p@a7vqV<;<:xTazy>aykRaR?vv2bA2mbd<n:8,D9VaQ-4qLqJ:j0O=7uQ7>i@h5xbuYa:szx0b|b?=E\\\"\\\",2):f(\\\"\\\"}>0gbhbXa7b\\\"\\\",2):f(\\\"\\\"}/n9QaYi3bV,Idn=S7B?w*+,bbO\\\"\\\",2):f(\\\"\\\"{Z:JwnzP6f8bb6bq2/*Oabbr*qqfbd,y\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}b667vfbFal9jblb<s6bYrbb4birM=6b8p1\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{btbOaz>8bOakui:>a3sPae;TaH9*>I\\\"\\\",2):f(\\\"\\\"{DqVakbUa|bD\\\"\\\",2):f(\\\"\\\"{FaH4XaOaY\\\"\\\",2):f(\\\"\\\"{avd*w871A<0b<a\\\"\\\",2):f(\\\"\\\"}oXa5bibJ+JyduGm4pUa\\\"\\\",2):f(\\\"\\\"}b?wybjb=p5bR6x9e;BuW5X,\\\"\\\",2):f(\\\"\\\"}uki\\\"\\\",2):f(\\\"\\\"}*x*k1998.-9-bwbdb"));
$write("%s",("kbx|G=mbmh>9hb@aBwfb4b*5j/6bSz3b8bubn\\\"\\\",2):f(\\\"\\\"}cb<tGgSz*uQa56>ajs5pI<Mol=Sk|bgq1zEaub:w3bZ|wbLyXs:\\\"\\\",2):f(\\\"\\\"{q|+60bOz2hX1KrIr\\\"\\\",2):f(\\\"\\\"{=32Yao,c2wbzoybb/Fa5b9/xb\\\"\\\",2):f(\\\"\\\"{bb/N<0b*wkblbo;y\\\"\\\",2):f(\\\"\\\"}HwOjUpTakbbbKwsr8b=aFa32;wRakbur3b*bcbtbrv@a..mbx<QaN<kiWqgrC|-8Waa.Z,Aa3wy<P.xoAaVaOzvbAoTa|+|bRa28*ravN3n6L,e*=:0./yrsTa=aWadzvq0rX-ibHu38csWaTa@aiz0r|<7y28BambQ-PaWa@aSaEa/bjoibOaXaAo3bit-bvb=oDs7b*bz*awS\\\"\\\",2):f(\\\"\\\"}@rZa0+a\\\"\\\",2):f(\\\"\\\"{vb6\\\"\\\",2):f(\\\"\\\"}a4Ui7z/;lb8vcu<2\\\"\\\",2):f(\\\"\\\"{b7b>;P6J/wbMsgx0yx|K-e-Etn3N\\\"\\\",2):f(\\\"\\\"{5bjd>al:fg86kb?,?a0bwb\\\"\\\",2):f(\\\"\\\"{bUaV,9*9bAocbPa?aOt40Ew?0IzV5|:H-mbx|DtOaZ,nzS,cb|8Va8bWakuXyWa3-Bu8->+\\\"\\\",2):f(\\\"\\\"{bw9tbo3t9*\\\"\\\",2):f(\\\"\\\"}7|W3Mw,b=aex-b7bKuP9Naz--/1:wbEzy*4bfb:x\\\"\\\",2):f(\\\"\\\"}b70jbU"));
$write("%s",("i8bFxibibi6j6::k6F,t8.7xb\\\"\\\",2):f(\\\"\\\"}bxvz-YaCacbkb9\\\"\\\",2):f(\\\"\\\"}*pXafb*b4bNa0b,bnojb8sW.zx\\\"\\\",2):f(\\\"\\\"}bjbX|W.OaybZa:txbL-Pa2bNakbxbZ4<*R|**\\\"\\\",2):f(\\\"\\\"{4Gaj5ZrOhOaWavb9|x\\\"\\\",2):f(\\\"\\\"{tbRaD\\\"\\\",2):f(\\\"\\\"}BazbXaIr28G\\\"\\\",2):f(\\\"\\\"{s.9-.dbbgvFavbk7Daibg\\\"\\\",2):f(\\\"\\\"}cb\\\"\\\",2):f(\\\"\\\"{bBaebUr>aHtwbh-0bCa06Ta*wo,ibWrZa*bxb.bQrZaxy1\\\"\\\",2):f(\\\"\\\"}Oa\\\"\\\",2):f(\\\"\\\"{bwb7bB\\\"\\\",2):f(\\\"\\\"}l2fgAu2w9bj+23=ajmUaDuPa.b;rOz<87pabOaPa=aDaXa1bkb;r|b5.kb5b98fb7bB8ubwkW-ZaebAoBaGaZ*hpP2vbYa6-+bmot\\\"\\\",2):f(\\\"\\\"}8bFa0bDao+n3@1Ca3bVaTay./baqiqlbDt\\\"\\\",2):f(\\\"\\\"{blzXatbx|46avIxu/w/61M3>o/b;6C\\\"\\\",2):f(\\\"\\\"}ohkiV/,b2b@fAiyk8b3bzbL7uqibf7vbr.fboh32*2M7bb8b\\\"\\\",2):f(\\\"\\\"{bgb1b1p9bU1moVz;5lqQrz0>aabutz4hv.7*\\\"\\\",2):f(\\\"\\\"}@fwbh+CrizSqwbH6yb.bj3.b@azz6b=sbbib4bCwF.ki:5?a"));
$write("%s",("vbabV6ykUaU1Tsfwn1@hCwb7C-1b<aUaz,RadzVzT3xrH6QawbabmjSavbgb0bFiZskr<aU1cbp*s||1Ta\\\"\\\",2):f(\\\"\\\"{b8bP\\\"\\\",2):f(\\\"\\\"{FaBf7ulqu10zrqbbBaxbGvL2\\\"\\\",2):f(\\\"\\\"}b06hb?0zb|bx|Wa7uzo.bZsQa<alqNax|7beqVa<tV5gbT5R5ZaP5Z,Uq\\\"\\\",2):f(\\\"\\\"{to\\\"\\\",2):f(\\\"\\\"}yb=lJ3g*=lH,L,M,K3K,f*t/,bJ1Axy+0xn\\\"\\\",2):f(\\\"\\\"}>v6bXaTaVni1Va5|G5Aalb.oub.xhbgsL\\\"\\\",2):f(\\\"\\\"}Kulb8b2wAo8bzy+04,so73Bu,oAo5bdwYaOzEaybxbAfcwTaCac2,b=pC\\\"\\\",2):f(\\\"\\\"}8vXajqHgJydbFx0w2,zbcbh5fbXaB+Wa2b8bn\\\"\\\",2):f(\\\"\\\"}T\\\"\\\",2):f(\\\"\\\"{kiO1fcZaablbR|WaCr;rv\\\"\\\",2):f(\\\"\\\"{/bwbP+aohbhbq1Xa=aZ-x+=a,bRabpOaQa432bki.46bEaebRaKw:-4b5b9,-d\\\"\\\",2):f(\\\"\\\"}b4bE32jbbWaMrkbSu6bs\\\"\\\",2):f(\\\"\\\"}7kAo<autdu@a2bYilbBfPazbmb3bD3+bZ2Qa0b,d-bDcdbVaJ.UaUaib4-\\\"\\\",2):f(\\\"\\\"}b.*Ec\\\"\\\",2):f(\\\"\\\"}xabYa4b,b=oHrebOo1bAon*?adbq.vn\\\"\\\",2):f(\\"));
$write("%s",("\"\\\"{iI3tn51Nx81eo<a*b@p2baidbldgu7k+o+rTaC|3zFgibCaQa8b6b-bkbSc@p7kjbKt=ahbx|jbauzbtvo*F1fb8b>aH-*bmbCaeb8b/b3\\\"\\\",2):f(\\\"\\\"}2v\\\"\\\",2):f(\\\"\\\"{tvb-0dk\\\"\\\",2):f(\\\"\\\"}u-wSsAoj,H2F2Qa9b.bZn*b2bKr<a2b@hybZpwbRn.blbj,BaKz*bkb|fj/v*k-RazbP|\\\"\\\",2):f(\\\"\\\"{b?+lb\\\"\\\",2):f(\\\"\\\"{u/bkzpq/b\\\"\\\",2):f(\\\"\\\"{b<0kb2b\\\"\\\",2):f(\\\"\\\"}bSaAalokpY,W,0bNa0re-gbTaUy-p>oY*7tg-ZbZn7bjplb<yg2+bBa/be-c\\\"\\\",2):f(\\\"\\\"}8b\\\"\\\",2):f(\\\"\\\"}urwY1jbubAt\\\"\\\",2):f(\\\"\\\"}qsl*b.bbbtbSzibkiK1Ao\\\"\\\",2):f(\\\"\\\"{b2bvuAsAaubXaFa*tCa+bwb+yPa\\\"\\\",2):f(\\\"\\\"{bfbEa?pkb,b<\\\"\\\",2):f(\\\"\\\"{3\\\"\\\",2):f(\\\"\\\"{h*41.\\\"\\\",2):f(\\\"\\\"{rnI,x/ZaCwfb5g9*S|7bfbabUu2b<akbYa@hQxj*BaabFvjbPa3beb:v@ax\\\"\\\",2):f(\\\"\\\"{ybYa60+bFv1brrSa<aFawb2bab+b8.rujxOjFvTa+burzbj*GaG*+b:r7|dlCav*hoab+dhzDaohx|wbkbwq@aqoV|B\\\"\\\",2):f(\\\"\\\"}tb>a1bYa.bn\\"));
$write("%s",("\"\\\",2):f(\\\"\\\"}bbi\\\"\\\",2):f(\\\"\\\"}Qx|bOa1b3\\\"\\\",2):f(\\\"\\\"}Ca.xDi4y*b/bYrQsA+SahbjbAo3phbAohc3yYv2bjbgbg05.N/c0K/Qa>aY/Y|L/kiS/T/Na>aQ/SaL/AoAoL/5b?/\\\"\\\",2):f(\\\"\\\"{bcbgbjwwbAowx-blbCq,.j/0.>a1htb-o...bcb0.q/m/p/l/j/rs5b0bjbRa4bvbfw=a\\\"\\\",2):f(\\\"\\\"}.s/0.vnL,+\\\"\\\",2):f(\\\"\\\"{G,evC,GxAop/qsr.Qa0.rs0.OaEa.b-.<y7b+b1hFyOaW,ybOa0.?ayk?qDaZ,<aWaI-?pBa1hBaF.>aG.E.@a7b5mW-Pn@a1b@ajrr.YaVa--r.,,/bVaPa>aEaq,=a1hRaVaUa?amb=aEaZ,bms.TaSa@agbNaSalbRa.bSadbxb.oOamb>aSa0hYa0bBa=agbUaEaSaWamb@aRaTsKtCa|zx+WaKtE|.b+zab7|.bRaab=oZrNwabFadbVnjyl\\\"\\\",2):f(\\\"\\\"};w=y0bxqOafbZa1bib?a\\\"\\\",2):f(\\\"\\\"}b?aCyT||bxbRa6bstxb6bNa@aQa6b*bboBa\\\"\\\",2):f(\\\"\\\"{bbbSaTaOalbxuPaVa\\\"\\\",2):f(\\\"\\\"}vOaYa<\\\"\\\",2):f(\\\"\\\"{/bZa4bkb3b+qibWalbgbN\\\"\\\",2):f(\\\"\\\"{lbPa7bDtn+hbUaOaXz,b3\\\"\\\",2):f(\\\"\\\"{4\\\"\\\",2):f(\\\""));
$write("%s",("\\\"{E,c*onMx/\\\"\\\",2):f(\\\"\\\"{3\\\"\\\",2):f(\\\"\\\"{-\\\"\\\",2):f(\\\"\\\"{0\\\"\\\",2):f(\\\"\\\"{2\\\"\\\",2):f(\\\"\\\"{b*jcXzL\\\"\\\",2):f(\\\"\\\"{wk7,2b*bTs-b*bjbOa,bzbYa/rebEabbUa7bW+wblb6b6bvb>owbQaDw+bftPaebUaAaOadbQaPqtb*bzb/bRaUa0b?a/\\\"\\\",2):f(\\\"\\\"}abxyjtxjQa7bcbRa9b,bOrzbNa>x\\\"\\\",2):f(\\\"\\\"{bxvSa4bhbWaUa8b,jVa4bDa2w.txb=a\\\"\\\",2):f(\\\"\\\"}b/b@avbX*P\\\"\\\",2):f(\\\"\\\"}N\\\"\\\",2):f(\\\"\\\"}ubUa4bYaDaubWatbnuSaeb6bwb9\\\"\\\",2):f(\\\"\\\"}PaTaAazy\\\"\\\",2):f(\\\"\\\"}bbbRa@ahbFa9blbJsk+,b.*NazbZaUaPa1blbUaRx6bOaAo+bdbR\\\"\\\",2):f(\\\"\\\"}R*:wAoOy-bOz;kAo0bv\\\"\\\",2):f(\\\"\\\"{Oa3bbxfbvb<a1bVqR\\\"\\\",2):f(\\\"\\\"}Ttibzbub?a.btbMw0b/bubmbfwdw0b+bjb1h6bjbeb2bPatblbkbcsgpW|AolbpjcblbmbbbFakbItLh7bQadqfb\\\"\\\",2):f(\\\"\\\"}bvbibYhslAaav>lLx3\\\"\\\",2):f(\\\"\\\"{Jx3\\\"\\\",2):f(\\\"\\\"{|sKxucN|qzbb\\\"\\\",2):f(\\\"\\\"}babCavb=aki@oyb\\\"\\\",2):f(\\\"\\\"}by\\\"\\"));
$write("%s",("\",2):f(\\\"\\\"}/bCaI\\\"\\\",2):f(\\\"\\\"}1h0b0w*uRa8bhbtbeb\\\"\\\",2):f(\\\"\\\"{v9byb,bAw?wcbAa,b\\\"\\\",2):f(\\\"\\\"}bQsnzVpYakbib<aebkb8bBaXa;i/bvb;zCa0bZaAafo:w/bDaebzu5pjb7bBavbOaIq-b=aIrZazb4bCaNaqxUaAoOaxbmbmbZt5bmbybNa?aFa*b\\\"\\\",2):f(\\\"\\\"}oQattXa2bks7oxujbTaUaabEaJ\\\"\\\",2):f(\\\"\\\"{dbUa\\\"\\\",2):f(\\\"\\\"{b+d5b-bJoXaZahcTa8guf7tDaPaY2db+|Ca4u5b;wvbsq?ab|abtbN\\\"\\\",2):f(\\\"\\\"{ab6b4b>xFaOa\\\"\\\",2):f(\\\"\\\"{v.bPqeb|bmb7qbb/bkbfu|ydbib?zpw>a+blbEavbqo\\\"\\\",2):f(\\\"\\\"}bib@p\\\"\\\",2):f(\\\"\\\"{b>aYabb,bOa@pzbAoCaWaOa9pdb,bRvNy7gVo9bZa>aZaBa6\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"}b|rSaavbv,\\\"\\\",2):f(\\\"\\\"{Zu\\\"\\\",2):f(\\\"\\\"{sOxysav*szsHx-bjbYix\\\"\\\",2):f(\\\"\\\"{NaegUalb-bAuBawbwbUaPulbYzWz,bb\\\"\\\",2):f(\\\"\\\"{GaVx+bvbgqQpmtZa6bubNa+b*bib5bNa-bEawbNaOa0b/z-bJw9bub3buo4b1pPa\\\"\\\",2):f(\\\"\\\"}bAoeg;xYaub9oybyb+b*v<atba"));
$write("%s",("b8bDaKh?afbibwbXaRauyZplbebEw.bvkgb2bAa8yizHq4bXaSacbCyQq7bdbabTa3bubPaurXasqOa/bNyVaku/bAambwqlbXaybkbAa.bDaNa2bBa.b8bYxzbRa0bxvOa>a?a|b=a\\\"\\\",2):f(\\\"\\\"{b*o3bCaAo2bpxPwOaOr<smbkiktAaTaebJt9bfumb1bsrEambgbhqBaWakbZa5bDt*bSsib.b>x,bWa1bcb3bykbb1b?axtVv4bdbqx>xSxaxkv?vDtNaYaZa\\\"\\\",2):f(\\\"\\\"{ixpypyiwpavcvavdv.bBaxj9bBa>xtbBatbgb/b8vPa6b8bjb:q=oPaub7bTaabkbbuebhc<oxx6b,bVvdb0bAo*bRaBa5b8bEiHqAatb9b\\\"\\\",2):f(\\\"\\\"}b3bHt/bOaubgbmb/b\\\"\\\",2):f(\\\"\\\"}bgbTr-bkiUwlt\\\"\\\",2):f(\\\"\\\"}b2bGrNs|rufZaQu=abb0bcb5bYafbQa?aIqwbSaBaFahb0b3blb5b=aCadb=aUtab2g:i8bEaWaVa\\\"\\\",2):f(\\\"\\\"{bPa\\\"\\\",2):f(\\\"\\\"{txbEa0b,vBa:p7b\\\"\\\",2):f(\\\"\\\"{bYa\\\"\\\",2):f(\\\"\\\"}bdbyb/bfbPa@a|babhbVqebslDr,b7b3bBa0bRaiblbxbib>aAo|bjsdb5bZa9rhvgp<aubjbab7bvoPakbgvcbvblbQotbNaBa+r\\\"\\\",2):f(\\\"\\\"{b-b5bybYoabcb7bXaQa"));
$write("%s",("gpAqdb.bWaYa,b*bTaVrOaTutb\\\"\\\",2):f(\\\"\\\"{b/bcb6bmbBagb5bOaCa=a+b5bTa<sOa|bAo-bBq@q/bUaavwsYuxs4a\\\"\\\",2):f(\\\"\\\"}s<luscb<a\\\"\\\",2):f(\\\"\\\"}bYaQa\\\"\\\",2):f(\\\"\\\"}bIgbbDaFovbsr6bZajtku|b,qXa/lxbeb5bEa>p8bFs*bEaCayb8bhhRaBfjpYaHrdb0gWaooPaXa6bibmbxbgbkbWaRa5bdrFaUaUnFacb1b7bxj8bebXaDa2bmbXacb8bZr9bmb0bkbSa4t\\\"\\\",2):f(\\\"\\\"{bDt7bAoeb2gdtmbEjSaSaXiVaSa3bYacbibPoab\\\"\\\",2):f(\\\"\\\"}b+b/l@aAa3bPa|b6bkbFa?a/b-bRaSabbwbRoPoWa8b7b4bFgEiRaujXaabwbAfVapqnq7bNa.b<r.l/b7bEa-bAombwb1b2bCo+buo@aXavb\\\"\\\",2):f(\\\"\\\"}bzbeq7bSakb3sOaab,d6b.p-b\\\"\\\",2):f(\\\"\\\"{bubfbzb@aBa>aGqEqXa+bGiibAoYaeb.bab4bPaxbFa/bPaJd+bFa>a8p5r3rSa8b0r.rvnyiupvsvpzptpvnvnMinp,r*rUaVa5bRaXa.bLpib6bSafbbbQaUaPnabzbWaXabbBpbbcb\\\"\\\",2):f(\\\"\\\"}b@acb1hvbjbcbUa,bTaNa5b3b,bAoyoYaFa|bNqub8b-b9bPa+bTa1bFa.b8pebyo1bfbSqUaQa."));
$write("%s",("bibhbQa\\\"\\\",2):f(\\\"\\\"{b.b?aab<a9bvbzb@qTaYa-bmb\\\"\\\",2):f(\\\"\\\"{b4b7b8b2bfb-b3bUaki:oVa@a*bwbvoQaybDa@aAoPaibdb2h8b?a3b>aibRa/bWa\\\"\\\",2):f(\\\"\\\"}b1bdb8b.bTaQambebebQa|b\\\"\\\",2):f(\\\"\\\"{bkbxq/pNa\\\"\\\",2):f(\\\"\\\"}b5b@aFa+bEaEaFaaqYp>oYi5bDa1bub|bVadbao\\\"\\\",2):f(\\\"\\\"{bLogb4bjbNaNhkbRavbdbublbvbRa\\\"\\\",2):f(\\\"\\\"{bebmbibTaGpFagblbVacbYaabNaTo|bhb*bBaDajbtccbTa-ptbCatb2bdbTatbDaDa3bAa0bdbCa>aTa8bNa|bAaFa4bBfbb|b*bDakb4b>a,bZahbDaxbcb?a\\\"\\\",2):f(\\\"\\\"{ippqp8lop8lrpun\\\"\\\",2):f(\\\"\\\"{iynzn\\\"\\\",2):f(\\\"\\\"{ixnvn9f-htbdbZakbebZa,bvbcb+bfb.bmbtb|bBajbjb\\\"\\\",2):f(\\\"\\\"}bwbEa1bebegkbdbkdEa9bwb*bYa7b|blbGa;ogbvbNa1bkiqb7b<a>adbBalb,bYa.o/o-o+o7b/bYagbibjbDavbDaQaEa+d0bybgb.b-beblbzb,bNa7bvbCaEahb<aCabb*b8hQaub*bWaQagbSa,bEa7b6bAaEaXlBn1nJm\\\"\\\",2):f(\\\"\\\"{mym*nXfMm-m<n;afn.m?a,mfnLmJl"));
$write("%s",("6n-bXlCmCaIlcnwbicfnKlxm-nEaimMmzmIl3mumsmvn@l@lpn4asn9ayiqn8lnn;l\\\"\\\",2):f(\\\"\\\"{i?l/b\\\"\\\",2):f(\\\"\\\"{f-a;hub@h8aDmQm4mVmHl9aEaOaMmKm<m2i:a-bMm=aAa-a=m7mCaimmm2m@a<a-b|e@m6mamwmlmcmamYl*m5m:aCa|e/m>aAaxmhmcm9aFldmAa:kTl|evm/lXlkmBa-aZlSlQl*bvbtb/b-a+bIdLlemMlVl@aTlXlSe|eRlWl?aAaIl\\\"\\\",2):f(\\\"\\\"{bGlNlLlFaJlHlFlHaDl9a|eElxb8a+e-a1beg8aXf,l8arb|eidxi=l=l9l3aLiyi7l-fziylOhFf6b-a+czbxbubHaqb6aqbEiFiDi5aqb@g-a,bAfzb.bKfnbxb\\\"\\\",2):f(\\\"\\\"}ikiZgXg\\\"\\\",2):f(\\\"\\\"{gag\\\"\\\",2):f(\\\"\\\"}h6hjk7jqk?a=aLi;dLfbk7i?kvh=ktcBa3aPhIgDiwbPf?a@krkWjBa?aKi6e;hrbck7hDhZj*hXjDa?a>aKi2b3bGiUfyj8f2i-bCjCa3aKa\\\"\\\",2):f(\\\"\\\"{b;a3gwbccIa3b1b-j,b|b0avhakik5jCaKi.bti7hvhQiOiMi@aKiyb3bTj?a9j5i5h6jBaLiMf1i\\\"\\\",2):f(\\\"\\\"{g\\\"\\\",2):f(\\\"\\\"{gsbubwbki-aDjBj:a;b?j1b0b-b3aAa3a7b-aki.a:b:b,b7hWhPimiNi@"));
$write("%s",("a3a;hwb+b-aPcuj/b8b1bPcxb;aUf-b:fZapg|b.b5b-amj>i3bWfvb|bIgGipgfg3bgf;a<b:b3b-a8bIg,bxb2b2btb;a7h*h6iPa4i3a>a3a5anb-aEi/b3b4b.bHa8byb2b2gtbWfxb5b+bYg7h5hliYhWh;d+cKfHa-i-iFaGaji|fld4a.gwi/auh4a-afgdgMaFa=aWh-bYhDhChGa+bJdRh9a/b5a|fCc8g-bPaBaobDhHfMa9aMaIa5axb3b.b4b0bxbzb-btbeg7hkg5hGaMbHg2bzb;azbLfccJa7b?a?auh*hCdYaOaVafbVaibNa=avhvh?a;aSgVaNaUa.guhkgvbpbEa*c7bAaAa>aDa>anbJdubSczbPfIcQgyfwfuf2bsfNd3bHa?e-a-fZf:aIa+c9f:avbldub4bcb-b3ggc0gHaebdbJaGagfef8a1bxbwbtbxbUaac|b3bdgfb/akgzgtbxcRf?a1akg-a6a5bhg>azd:a,cNah\\\\\\\"\\\"),\\\\n(\\\\\\\"\\\"gwb.b;b>aagob,c:a-a.b\\\"\\\",2):f(\\\"\\\"{bvbxb5a1aob,fCe2b-a:b1dtbHa6a/c2b/a,fPcFf/b:b6aKa6e1b4eIa8btb1b1bNaGatb5a+ctb,b-a\\\"\\\",2):f(\\\"\\\"{fyb3dMd-aDdBd@dmf/aob5a.d,d*d-b4b7eSc;axb+b.bbcZb0cbfJasdHa/aed+e0cGb/d,btb-b4aWbudpcgdLc=chchd6are"));
$write("%s",("Oapc0cNb/a;bje/eGaHb5dedOb.a8aNd8aLdLa=a>aIaOaJapb6a+e5azb+cdcfbhc;aOaFdYd6aHaCa@aIaQd8aHa=a.cIbCbMd\\\"\\\",2):f(\\\"\\\"{cycvcocRapcXbocTa;b;bpbgbYdJaGbRanbQaJagbnbcb>dqc5dpbebnbOa8a0c4aJaTa5a+btb5bxbJaQa,c*cRa5a1bzc6aedMa0c3bldjd;aeded8ard5a6a5aedxb/btbvb2bxb,c1b4b3bxb1b0cocPa8aNapcMagdUc3b|b+b/b2b4arcFbnc4a=a?axbtc4aSbJcPbKckcic+bZb3b-bzcXbqcFb5aMa/ancvc+b+b|byb4a9cVbNa5aRb7cFbnbFbMapb2c.aMaFb.a4a5aJaOa-a-b|b-aeb5aicybHa<b/akc>a>aXb6aOb/a8a6a/apb4a1b.b3bvb4b1b3b2b-b.bvb4anb/aJaPa5a8a4a6apbEb5a5aB,ab,b9a4apbpbnb8anb4aGa=a:bJacb!\\\"\\\",2):f(\\\"\\\"})46(f\\\"\\\",2):f(\\\"\\\"{#~[2xha=s,y=z,13&X3^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\"));
$write("%s",("\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'yay,]99999[gnirtS wen=][c n3aea\\\"\\\",2):f(\\\"\\\"{)v]y3b&a(niam diov citats cilbup\\\"\\\",2):f(\\\"\\\"{RQ ssalcz4rfa cdlnl3c/a;maertStnirP/oi/avajL tuo/metsyS/gnal/avajm4bdateg@3doa2 kcats timil.v3dga]; V);Q4aC3ecaL[b5aX4hha dohtem?3e;4nga repus&3ecaRQ@3cgassalc.<5joa(=:s;0=:c=:i;)|4ajaerudecorp/3fqa(tnirp.biL.oken\\\"\\\",2):f(\\\"\\\"{.3bianoitcnufR6\\\"\\\",2):f(\\\"\\\"{sa(rtStup=niam^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^32^[2fha\\\"\\\",2):f(\\\"\\\"})3(f\\\"\\\",2):f(\\\"\\\"{#v3m"));
$write("%s",("ja13(f\\\"\\\",2):f(\\\"\\\"{#,4353(ga36(f\\\"\\\",2):f(\\\"\\\"{#j4[j4boa(etirw.z;)tuo.N8aba(67b~auptuOPIZG.piz.litu.avaj wen=zG4Zka91361(f\\\"\\\",2):f(\\\"\\\"{#tm4[m4c5aR0Z0Z/512152353/2/2166263=4/3141726??:1518191:1/@4[@4cda*6 Q5[p4dea1312^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'5[w8[$5ofa41310r4[r4c7=[B>[j4[^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'6pma(amirpmi oicy4[(5[j4hma++]371[]591[?6[?6cpani;RQ omtirogla\\\"\\\","));
$write("%s",("2):f(\\\"\\\"{4[\\\"\\\",2):f(\\\"\\\"{4cua;t:\\\"\\\",2):f(\\\"\\\"}%%%%\\\"\\\",2):f(\\\"\\\"}fi\\\"\\\",2):f(\\\"\\\"}*-84\\\"\\\",2):f(\\\"\\\"})48z3b(a]i[\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"}+17\\\"\\\",2):f(\\\"\\\"{<84.;i:-i602\\\"\\\",2):f(\\\"\\\"{;i:911\\\"\\\",2):f(\\\"\\\"{;j:632N4Zsa7218(f\\\"\\\",2):f(\\\"\\\"{#(tnirP.tmfIIcfacnuf;&4[&4bdatmfn4[n4cgaropmi;ILagagakcap~4Zea1304T6dbapD6[r4cba-l4[l4bjatnirp tesY>[ca89&AafantnirK7[ia959(f\\\"\\\",2):f(\\\"\\\"{#fp4[ga^64^\\\"\\\",2):f(\\\"\\\"})74[8awa,s(llAetirW;)(resUtxeT:Paca=:R6[ba1Q6ak8ap4[p4adaS Cn4[vEaca&(z5[z5aba 06[06[06piaRQ margo^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'5[t4cjaS D : ; R-5[%L[j4[j4o%6[k4a"));
$write("%s",("qa. EPYT B C : ; Az4[56[j4[j4nka)*,*(ETIRW/6[J7chaA B : ;s4[s4aba [2cr4[*5dia: ^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"' ohce4B[ka3(f\\\"\\\",2):f(\\\"\\\"{#(stup;Rcdatniy4/ca0153.ea%%%%m4[m4[53ipaparwyyon noitpoz4023[230ca(nVO.ba5FQa\\\"\\\",2):f(\\\"\\\"{aetirwf:oin\\\"\\\",2):f(\\\"\\\"})8(f\\\"\\\",2):f(\\\"\\\"{#>-)_(niamp3c\\\"\\\",2):f(\\\"\\\"{P)ka(f\\\"\\\",2):f(\\\"\\\"{# cnirp/L)l;eja.OI[p]^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^1"));
$write("%s",("^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'[(3rba@~Wa7;alaM dohtem06x*3c|5aV;cpadiov;oidts.dts &Ya;6n+4d\\\"\\\",2):f(\\\"\\\"{3kkaenil-etirw~5dva(,^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'s%^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\"));
$write("%s",("\"\\\"'(gol.elosnoc;)^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'73g\\\"\\\",2):f(\\\"\\\"}a^129^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"' nioj.)1+n(yarrA>-)n(=fI3cwa^31^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",2):f(\\\"\\\"}54,1\\\"\\\",2):f(\\\"\\\"{.^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"# qes-er()|3cH3bba^31^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\"));
$write("%s",("\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"p3lg3fw3hla1% ecalper.j4dea^128^+Ac/arts(# pam(]YALPSID^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\".NOISIVID ERUDECORPA3cma.RQ .DI-MARGv3g53d|bNOITACIFITNEDI^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"[tac-yzal(s[qesod(^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"))System.Console.Write($^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\""));
$write("%s",("\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"Put caffeine \\\"\\\",2):f(\\\"\\\"{(int)c\\\"\\\",2):f(\\\"\\\"} into the mixing bowl.^64^n^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");M3pva^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"Liquify contents ofE3oeaPour^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'3w^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'4e\\\"\\\",2):"));
$write("%s",("f(\\\"\\\"{abaking dish.^64^n^64^nServes 164cma\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}^31^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");\\\"\\\",2):f(\\\"\\\"}/****/e3a^15^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"),s[999999],*q=s;int main()\\\"\\\",2):f(\\\"\\\"{int n,m;for(;*p;)\\\"\\\",2):f(\\\"\\\"{n=(*p-5)%92+(p[1]-5)%92*87;p+=2;if(n>3999)for(m=(*p++-5)%92+6;m--;q++)*q=q[4000-n];else for(;n--;)*q++=*p++;\\\"\\\",2):f(\\\"\\\"}puts(s);return 0;\\\"\\\",2):f(\\\"\\\"}^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"))\\\"\\\",2):f(\\\"\\\"{s+=^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"00g,^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9"));
$write("%s",("):f(\\\"\\\"\\\\\\\"\\\";for(m=1;m<256;m*=2)s+=^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"00g,4,:^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"+(c/m%2>0?^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"4+^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\":^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")+^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\",^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";f(s);s=^7^\\\"\\\",57):f(\\\"\\"));
$write("%s",("\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"4,:,^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";\\\"\\\",2):f(\\\"\\\"}f(s+s);for(c:Base64.getDecoder().decode(^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"kaAREREX/I0ALn3n5ef6l/Pz8+fnz58/BOf5/7/hEX/OZzM5mCX/OczmZzBPn5+X/OczMznBL/nM5mZzBPu++fPPOc5zngnnOZzOZgnBMGAW7A==^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"))\\\"\\\",2):f(\\\"\\\"{c=c<0?256+c:c;for(i=0;i++<3;c/=8)f(c%8);f(^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"8*+8*+,^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");\\\"\\\",2):f(\\\"\\\"}f(^7^\\\"\\\",57):f(\\"));
$write("%s",("\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"@^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");^1^\\\"\\\",4):f(\\\"\\\"'|sed -e^1^\\\"\\\",4):f(\\\"\\\"'s/^16^/^32^/g^1^\\\"\\\",4):f(\\\"\\\"' -e^1^\\\"\\\",4):f(\\\"\\\"'s/^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"/^16^q/g^1^\\\"\\\",4):f(\\\"\\\"' -e^1^\\\"\\\",4):f(\\\"\\\"'s/.*/print ^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^8^nquit/^1^\\\"\\\",4):f(\\\"\\\"'^3^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")\\\"\\\",2):f(\\\"\\\"}^1^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\"));
$write("%s",("\",9):f(\\\"\\\"\\\\\\\"\\\")\\\"\\\",4):f(\\\"\\\"');\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\").split(\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",64):f(\\\"\\\"^\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");for(int i=1;i<a.length;a[0]+=a[i+1],i+=2)\\\"\\\",2):f(\\\"\\\"{a[0]+=\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",89):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\".repeat(Integer.parseInt(a[i]));\\\"\\\",2):f(\\\"\\\"}System.out.print(a[0]);\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";FORiTO UPBtDO INTn:=ABSt[i];print(REPR(50+n%64)+c+REPR(50+n%8MOD8)+c+REPR(50+nMOD8)+b+\\\"\\\""));
$write("%s",(",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"J\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"+a)OD\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"while(!=(S:length)0)\\\"\\\",2):f(\\\"\\\"{\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans c(S:read)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"D(c:to-integer)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 35 39\\\"\\\",2):f(\\\"\\\"}\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 24 149\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"interp:library\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"afnix-sio\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\""));
$write("%s",(",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans o(afnix:sio:OutputTerm)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"o:write B\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");end;\\\"\\\",1):f(\\\"\\\"\\\\\\\"\\\")\\\"\\\",1):f(\\\"\\\"nsys.exit 0'}\\\\\\\"\\\")\\\"\\\",0)]]></xsl:template></xsl:stylesheet>\\\":s.WriteByte(Asc(c)):Next:End Sub:End Module\")\nput=s\nprint\nqa!"));
end endmodule