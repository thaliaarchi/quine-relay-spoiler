module QR;initial begin $write("%s",("let s=(\"Module QR:Sub Main():Dim s,n,i,c As Object:n=Chr(10):For Each c in\\\"<?xml version='1.0'?><?xml-stylesheet type='text/xsl'href='QR.xslt'?><xsl:stylesheet version='1.0' xmlns:xsl='http://www.w3.org/1999/XSL/Transform'><xsl:output method='text'/><xsl:template match='/'><![CDATA[sub f(s$,n)print(s$);:for i=1to n print(\\\"\\\"\\\\\\\\\\\"\\\");:next:end sub:f(\\\"\\\"write,format=\\\\\\\"\\\"%s%s%s%s%s\\\\\\\"\\\",\\\\n(\\\\\\\"\\\"\\\"\\\",2):f(\\\"\\\"write{-}{txt}{echo -E $'(\\\"\\\",1):f(\\\"\\\"\\\\\\\"\\\"with Ada.Text_Io;procedure qr is begin Ada.Text_Io.Put(\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans B(Buffer)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans O(n)\\\"\\\",2):f(\\\"\\\"{\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"B:add(Byte(+ 128 n))\\\"\\\",2):f(\\\"\\\"}\\\"\\\",9"));
$write("%s",("):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans f(v n)\\\"\\\",2):f(\\\"\\\"{\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"O(+(/ n 64)107)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"O(n:mod 64)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"O v\\\"\\\",2):f(\\\"\\\"}\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans D(n)\\\"\\\",2):f(\\\"\\\"{if(< n 4)\\\"\\\",2):f(\\\"\\\"{f(+(* 6 n)9)48\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{if(n:odd-p)\\\"\\\",2):f(\\\"\\\"{D(- n 3)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 27 48\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 36 11\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{D(/ n 2)\\\"\\\",9):f("));
$write("%s",("\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 21 48\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 48 20\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans S(Buffer\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"STRINGz:=REPR226+REPR153,a:=z+REPR166,b:=a+\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"2\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"+z+REPR160,c:=b+\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"8\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"+z+REPR165,t:=\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"#include<iostream>\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"+REPR(10)+\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"int\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"+REPR(32)"));
$write("%s",("+\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"main()\\\"\\\",2):f(\\\"\\\"{puts(\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"class QR\\\"\\\",2):f(\\\"\\\"{public static void main(String[]a)\\\"\\\",2):f(\\\"\\\"{a=(\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"write(\\\"\\\",4):f(\\\"\\\"'implement main0()=print(^1^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"BEGIN\\\"\\\",2):f(\\\"\\\"{print(^3^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"echo ^1^\\\"\\\",4):f(\\\"\\\"'f(s)\\\"\\\",2):f(\\\"\\\"{System.out.print(s);\\\"\\\",2):f(\\\"\\\"}s=^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"389**6+44*6+00p45*,^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9"));
$write("%s",("):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";for(c:(^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"#include<stdio.h>^8^nchar*p=(^15^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"Ra#include<iostream>^16^nint main()\\\"\\\",2):f(\\\"\\\"{std::cout<<(^31^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"class Program\\\"\\\",2):f(\\\"\\\"{public static void M83abbSystem.Console.Write(^63^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"Quine Relay Coffee.^64^n^64^nIngredients.^64^n^63^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");for(int i=9;i++<126;)[3pva$^63^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\""));
$write("%s",("\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",2):f(\\\"\\\"{i\\\"\\\",2):f(\\\"\\\"} g caffeine \\\"\\\",2):f(\\\"\\\"{i\\\"\\\",2):f(\\\"\\\"}I3b54rja^64^nMethodv4f#aeach(char c in(^63^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")))^127^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")^127^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^32^[2al3dp3c[2cs3c,3l[2k@3kqa^31^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")s rts(ecalper.h3eja^127^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"     53c4a SUTATS(egassem^127^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):"));
$write("%s",("f(\\\"\\\"\\\\\\\"\\\"rts(nltnirp(])]^127^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\".NUR POTSu4cba.C3dh3dX3bba[65bX4df5lp3lna\\\"\\\",2):f(\\\"\\\"})1(f\\\"\\\",2):f(\\\"\\\"{#\\\"\\\",2):f(\\\"\\\"};)06xt3dba;+3noa3(f\\\"\\\",2):f(\\\"\\\"{#qp]\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"};)0,#3rv3rR3sv3mba723284-fa(f;)1q5.ba.>4[ga#(f;)3P6[=43ba7=4.<4[<4[<4[v3gJ=d=4[73++>u?4[73xda,43?4[?43ma^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"' D ; EYB RCo8[.6[?4;ba5qB/daDNE&6[&6[&6[8Emca AL9[)6[)6[v3oeaPOTS^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\""));
$write("%s",("\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'6[^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'6[^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'6[M9pL9[(6[(6[v3moaRQ margorp dne16[16[16[v3lbaST9[&6[&6[JQ[~6[?4Nba4~6[~6[~6[~6>ba&g=[$6[$6[.@neaPOOL|N[,6[4@[>Xp>4[#6[#6[#6[#6[#6[#6\\\"\\\",2):f(\\\"\\\"}da&,)l=[^1^\\\"\\\",4):f(\\\"\\\"'^7^\\"));
$write("%s",("\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'6[^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'6[eUnga. TNUO9@[,6[,6[83nearahc1G[)6[)6[R9ogaB OD 0hU[-6[-6[%No33)$6[$6[%NBca)Av=[&6[&6[HQoCQ[^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'6[p=[v3nqaEUN"));
$write("%s",("ITNOC      0136[36[36[sDnV9[&6[&6[lDoG@[^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'68l41ba0l4.27[275gaS RC .47[X:[)6[@4mja1=I 01 OD-6[-6[-6[NAneaA PU*6[*6[*6[v3:~6[~6[:OBxa;TIUQ;)s(maertSesolC;))T4[96[?4:ca11Y9/fatiuqnq41ca82p;[57[57[?4jda932A4.172ca65m4/i<[27[gC<ba9D?/maetalpmetdne.>72da215>7[>7[>7[?4kca007?/ca\\\"\\\",2):f(\\\"\\\"};^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'6[^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\""));
$write("%s",(",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'6[?4<ba8A4/#X[j47da862E@/batX6[=8[?4:ca44OPY>8[cCkda283m4[x5[bDgca8757/%a315133A71/129@31916G21661421553/:9[\\\"\\\",2):f(\\\"\\\"{;[9M;ca99\\\"\\\",2):f(\\\"\\\"{;[b9[\\\"\\\",2):f(\\\"\\\"{;[x5[v9wca2357/ra%%%%\\\"\\\",2):f(\\\"\\\"}*+1%%%%811 -jX2ca84;D/;6[T8[x5[j4Fda688T8/haj:+1 j@w?[W@[?4:ca02W@[D8[b;[x5[b;xca0457/baww9[W:[?4:ca60ZB[>8[W:[x5[2?zl4WU:[U:[?4mda398U:[<8[U:[x5[57wca34l4.baWv9[V:[KX;ca73=8[=8[j4gda277x5/ba\\\"\\\",2):f(\\\"\\\"{Y6[>8[2P;c</<8[8@[x5[3XHba2x5/wa)(esolc.z;)][etyb sa)^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\""));
$write("%s",("\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'.9[o;[?4:ba5jT/#6[#6[#6[#6[#6[7GMba4TA[;?[TA[x5[x5[x5[x5[x5[x5[x5[x5[x5[x5[m4[x5[x5[x5[x5[x5[x5[x5[x5[x5[x5[x5[x5[m4[x5[j4cda267iT[iT[iT[-W[#6[#6[#6Rba,%6[%6[%6[E9[#6[#6[#6~ba!m41ba6m4/ca~~37[37[37[S:[#6[#6[#6~ea(rt.(6[(6[(6[H9[#6[#6[#6~ba)BA[v3cda\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"};p4[SBfdadnes4[s4gra~~~~PUEVIGESAELPnr3ala~~1,TUODAERw3a:4[:4i$a(etirw;\\\"\\\",2):f(\\\"\\\"};u=:c;))652%%%%)u-c((||54[54ida#-<u4[u4ida||i15[15lhaBUS1,ODz4[^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\"));
$write("%s",("\",4):f(\\\"\\\"'8pka)3/4%%%%i(g:c4;[04jr;[r;wPa2=:/t;2%%%%t+2*u=:u\\\"\\\",2):f(\\\"\\\"{od7 ot0 yreve;i-=:u;1=:+i\\\"\\\",2):f(\\\"\\\"{od))1(evom(dro=:t elihw?s;)s*z9[L;ny9[y9uz4[z4i0Adladohtem dne.s3dganrutern3dCaV);gnirtS/gnal/avajL(nltnirp/maertStnirP/oi/avaj lautrivekovniJ3d25[25i[2cib\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"};0=q;)]q[c=z(tnirp.tuo.metsyS;)0(tArahc.y+z=]++n[c;y:]q[c?n<q=y\\\"\\\",2):f(\\\"\\\"{)0>2%%%%++i(fi;48%%%%)31-)i>3c&as(+87*q=q\\\"\\\",2):f(\\\"\\\"{);23312<i;(rof;n)rahc(+O5[O5q[2k.4[.4%oa=]n[c);621<n++z6aqa0=q,0=n,0=i tni;R4[R4%oc6agi4asdRbQeclxfvfVk?f<bedPdoj\\\"\\\",2):f(\\\"\\\"}b;agb-a|dzdxd?fGb8aqeRdYd5a\\\"\\\",2):f(\\\"\\\"{b2b5i;agb-epb>aqeRdHa>aJaRaAdteFbae:b6aOa5aacsg+TaK9a6*4aLa7a;a4a<a=hcmkdxd;aNa?c6a|eebHaFaIaebzeJaeb9a/a6a2dQbUe-f2a-f9a6*5d6cRb"));
$write("%s",("C3gAc-f/aof0f?fSg7e\\\"\\\",2):f(\\\"\\\"}h4e.b2e6aRa;dSMVfz*5h;aTapc4aLcEegiof6amc6a-f;f:lsbdhIuDfybxcxc>aGaUeAa2a6ajg7a6a@ahg:a?aMbKaKa6a?e:aP,2aigGfMbIfTh>a:b1angamBf\\\"\\\",2):f(\\\"\\\"{bHauco0k-oH6@oHEc+sJaMa\\\"\\\",2):f(\\\"\\\"}bJaeLEc-bJaJaUa-bJaMdJa8bPr;aS|TaKaS|Ta8bTarj\\\"\\\",2):f(\\\"\\\"}bRTSaSaJ49bKaS|O|TaS|#3aoaJ4JSJaLaJaS|1|j4c\\\"\\\",2):f(\\\"\\\"{a8bJ44bJ4:b6@oH6@+brj\\\"\\\",2):f(\\\"\\\"}bJaHa\\\"\\\",2):f(\\\"\\\"{3acaJSk3a+aJaGUVa;a8bRt:aUa:aPrdi@f>fBl4a4psbsb2be3^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'madiDa-aIu*b-a>6asavWUe>avjhgKaKaigGf|6cgaHf?jRf$6esasbdh*b-a/bxcHa|f>ke3cZb\\\"\\\",2):f(\\\"\\\"}bhgXghgcg"));
$write("%s",("1ang\\\"\\\",2):f(\\\"\\\"{bHa>k?f-e:a:a\\\"\\\",2):f(\\\"\\\"}bHa?ahgJa\\\"\\\",2):f(\\\"\\\"}b5aAdte@a1angri>kxcpb7anb2b:bhg2f.j@dCf6aNjxcHaSfQfOfVj-aBfrifi?f-fng@f|f>kzeAgfiHaLj;a/a2h<bmhEh<apb/a2hEhnb4C7b:bhg/awh:fnglgFani|bi>1ba0h>.4a1aTh3b:bhgJa7bHa>kHaUeoiCe|bxc3b0a:bhgIa|bzeJa|p6b#aQbfi<b=a-a8m*c3bxdUe=a-a?aJ+9ai3ehb2bMa7aZg|bXgVgTgRg9apbYgWgUgSgKcdc4ijjEivuydzb7aEa|b*k|kMa8m*cEc,dJa>a2a:b6agjykMa?aJ+*i+cJh6a33k[axdtb+bvbyg/a2h=aXhRa7ICd7IkbuoyCXh1kDh7b5aLj?fwbjjUe2b5azgFi4b-bhcbsRjRjOu0c/bxd+h\\\"\\\",2):f(\\\"\\\"}hVi<@aea6a2bd@gqc0lsT6ayn2a5a*lqTjg3hQkovxjDhBhfnHa1dmd9h?f1k;kHa:e1k;k+l<b3bxd6a*h5k=hxlHSShxb\\\"\\\",2):f(\\\"\\\"{iacPa;aEiccOqpbubld1bZbyvnbWfbjZiQhVz\\\"\\\",2):f(\\\"\\\"{jGkchEkuj<b<b<b4j:b*j<b<b,c9j6j7b-b9j<vAg3bDduk;i9a7bwg-a5bZ|,c9j=a9a7bc3q3e13eca1j13ceaM<xkA3c/3gdaJb@m3"));
$write("%s",("fma=a8mEj9a7bl8u3amaShjkW\\\\\\\"\\\"),\\\\n(\\\\\\\"\\\"i4k,c9ji3a=a-aJdy@Ng,c9jsb?fTjPk:k:i2jCa:i6aTjPkQjuj6aHk0kHjOksk<bzeVDceaHajgK5cca,k53cIa:k8k3a6a<bShJipT2b2a2a+PNjJkriwbjj?f@a>anc:e7b5aDf=anbNjybnk5a,bJa6apBa^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'aubJa7b5aCgwbjjHa:e-b9a9b9aYjNjfg>am3a\\\"\\\",2):f(\\\"\\\"{a@a@aNjfg@a>a:a|b9a0b9a@a>aWCa=a>e|b>g9bJa0bNjfg-b9aYj9aZCJa9bNjnbJa6a|b5a,b?f:e-b*k1J-a[;a&a-lq@QWdi+Pfg8bAd5h-a+P@qbb-a+Pfg7s3hhb+PKc,iP*xd6a-b9a8b9a7bJcJaybymW:>aJa*c@dxc?b,bzo>aJa-b9lteUe@a>aMR5aDcf4:atcJaubKdvuVz,b4b-bDgR:aiaDkBkmd9h^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\""));
$write("%s",("\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'7gLfNkLkpb;awbjjnl-lq@6F63RW+RsT5FMYJdHdplvn7n3lHl3m\\\"\\\",2):f(\\\"\\\"{ntno.7nFlRaubhp?uct-0fQZxetg,\\\"\\\",2):f(\\\"\\\"}bDag,px8x7\\\"\\\",2):f(\\\"\\\"{BA.pEa\\\"\\\",2):f(\\\"\\\"}pTaShKTL2dbvbOaEvoIT*tbRaTsibCnnAHQkp8xItQntIM/9bQFhb=a/pDahbDarL1=Daty.tzXkdnwA?ibspvbDa8<rLMux2@aMwA|,dLpuTq@6F2D4Fn<NYC5>B6brIH*,1Q-WtS>Z0Ta\\\"\\\",2):f(\\\"\\\"}Cx0/bo+|bH,YA*Elbg<y\\\"\\\",2):f(\\\"\\\"}EPZaibW/kqtbEae+5b.BbbrNK/,b0Q\\\"\\\",2):f(\\\"\\\"}CXL2|y3v4W9tbyr/ytbtul9:\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"}o-8@rbbK-5JTaibwpT*sAM.zb6bd.uqMz2b0pU8@ai7;<Wazx-9rN,d,dC7+bbb;\\\"\\\",2):f(\\\"\\\"}b9F>\\\"\\\",2):f(\\\"\\\"{sdzUMy3P1a<,b9bfb@+z\\\"\\\",2):f(\\\"\\\"{hL"));
$write("%s",("GVxpq/s.Luuo/bW>9-K-jjeCYRQrr2RBl9\\\"\\\",2):f(\\\"\\\"{*EaHDI18*=5fWdS@|BQ*TY4b\\\"\\\",2):f(\\\"\\\"}*of=z<WaVasA,yv+8x-bf\\\"\\\",2):f(\\\"\\\"{?Kg,\\\"\\\",2):f(\\\"\\\"}C8,sAii28cvd.bbbJvnsFa.ii-qZ5@,u.KEaMI;pib+pUnacGn@BCy,kTa0bj5lbX>W/I<F\\\"\\\",2):f(\\\"\\\"}vWzPjb?aiy/.FP1uuw@ac.?2vq;NqFNv\\\"\\\",2):f(\\\"\\\"{zSae+W*ZX\\\"\\\",2):f(\\\"\\\"}o<oXawpcz-+FOdS9kTaAa,yGnQwJ,o+h,n/y@-bsr?rcy8JII*h@WB3Da8b\\\"\\\",2):f(\\\"\\\"}b5xJod6=GdQgUYa=GRSoxHnZXwbRag,vb-.FPDPHIW:APUsm0B3O.coaoA*DaPa6PYBEaT0j@UtTa@+Rag,@H2odrlbs6w6DaF/g,vb<oZzl1+H\\\"\\\",2):f(\\\"\\\"{tubY>Da~6e~dVao.hqEa8/nL5N@yMkOPF7:xmwX>/bYB\\\"\\\",2):f(\\\"\\\"}FDa|7QOubShxoDar6Daw6DavbS.HO<\\\"\\\",2):f(\\\"\\\"}DO4bSa2:28TsCvKCjb6mgbjbLo<26bCaR41Vgbjbvb>,xs7=Z,=aEabj\\\"\\\",2):f(\\\"\\\"{B\\\"\\\",2):f(\\\"\\\"{BE3CvTa76sQtOVa=aEaqOoOybfhqIZ|,XQxhO,bfOg,IClo@wjsl?eojDUNB3QaCveo?6QnNNg"));
$write("%s",(",ejTaJNSajb|NB36/Oag,f=QnoGKqKTNag,EqsVWn7Jlbvb5N+52N7L9bPa.N|NCn8b1tTazbn,iW8<b\\\"\\\",2):f(\\\"\\\"{n,ubz35s<Lsp*6eHbz3sv<LspgrAayCn,ubgrEa1bgb-|@aVa3bhbgN9bEausWv153\\\"\\\",2):f(\\\"\\\"{Ta3\\\"\\\",2):f(\\\"\\\"}?ahr,bACL2Y>-bo+Zz.rWplHyb7bw<zu?ehLX8z3oLZzRaubAakU*1qsf;:*DaNgzX;,h4OnPL,p6m=aPr?YPaDatbKpspyB5S,km3awaB<=aBT7pZzNkB<<ajbDS3o#3e~dDaHIA?Sp\\\"\\\",2):f(\\\"\\\"}AXLmu?pA9?pdb@?NkDaGnCao5ZaDiJz?aDaMxxbNn0bj*opTaPotbG8e|Y-+dip@a0qZaqQ/yo?,zv6JCT5<pEv:+Qo/i+P\\\"\\\",2):f(\\\"\\\"{Jq@QWXrhOG8xKDa\\\"\\\",2):f(\\\"\\\"{1SCPnkbC\\\"\\\",2):f(\\\"\\\"}jbQMT>AxShNthbT/\\\"\\\",2):f(\\\"\\\"{xyb=aM0RF@aA7JFKs0QDBrHuwhb0b6-xUDaT/Xaeb-bWL5ZbUp=,kWpfhp=,k0LPvuwRaMnW0+S*b9wmQ>N?p4j.yTAaqpo/bp/hb|1mxLrmxHTmE8x8bX01bx\\\"\\\",2):f(\\\"\\\"}9bfbbjUGv2Oa8Xt,OZ=Gy3ejb;M8xfbir57-bq|5bu7mtBGTa<ac5x6jDoQQvdzebdzz\\\"\\\",2):f(\\\"\\\"{@>"));
$write("%s",("UM||XB.*GpGLJCqoW|y3GaHYNa*ul\\\"\\\",2):f(\\\"\\\"{|qg1l+l\\\"\\\",2):f(\\\"\\\"{jbcrSpHHSyMuO9epdjtSrptVNuYfb;8A?S<e\\\"\\\",2):f(\\\"\\\"{>24vFR6mmPQ@CaHz7>SS:g-\\\"\\\",2):f(\\\"\\\"{Ng8z,09sNk-R8bBiC\\\"\\\",2):f(\\\"\\\"}f|+bibtoauYa3zWa-@zy\\\"\\\",2):f(\\\"\\\"}Xu7H*5bgfa,U32PBa0RWLTz<oZ,KY=j@a?*HqgcSsIN-+R\\\"\\\",2):f(\\\"\\\"{HsIpQ.-VEGoOG*F7Ur\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"{Jyw|ufkxbjFvmqqI0RlDpu6IAq\\\"\\\",2):f(\\\"\\\"},eb:8ShaO|r\\\"\\\",2):f(\\\"\\\"}:wt1biBNa8R@\\\"\\\",2):f(\\\"\\\"{BA.p=CU42PBa@rx,abp7dbJF1b0?lbA3wb\\\"\\\",2):f(\\\"\\\"{53Nyzb-e1\\\"\\\",2):f(\\\"\\\"}b2NJy*,1zShJOFA:.6Pyb*b:h<a\\\"\\\",2):f(\\\"\\\"{bx6e~dc3ShKTT>U>5Xo3JSLZOaC<;vNgubT>dt:8DBSP\\\"\\\",2):f(\\\"\\\"}*ibl+6vebMw5bg<sw.pGadR>|Is\\\"\\\",2):f(\\\"\\\"}w4qMvQBUPhbXN|bufn/uNiWl7qyXw.-ebOanuhbKu|I912b5bBaXaldybQtQaQww0EP:xD@=a9bwX9<VqdOGzr-|qc8ShaOZ7Ev*q.b;CF/ub0bgy;CELFsfNWaK"));
$write("%s",("H\\\"\\\",2):f(\\\"\\\"{VbbcbcLA\\\"\\\",2):f(\\\"\\\"{9+f/qDbbN*4s@q2N:P|17bibx0WqMk0?YQ2MM|ibabXH*+QTNavW3*h*SMZa1bFat+?asw?q2rq4IRF9yuTa>\\\"\\\",2):f(\\\"\\\"}8**6e%aNaybZa5x\\\"\\\",2):f(\\\"\\\"}00*cUU|G*n4Axg4/x*t5*Nas3gMc5*xC7=0?4*AP@>27+XAqzbR.Uas2l3eb:oS5Saq|tbqFwpQwtl?*Za9bG+ebShaOtbR5yb6v1btb0bNaWrAF?a*:+bjb21ws\\\"\\\",2):f(\\\"\\\"{KAxxDSa.KHIK1HI.K5bRaF75q15wRJ+s5IrtzP*N*Nx5bEV,b2iFaZ/3bghyb5b\\\"\\\",2):f(\\\"\\\"}47|Ta,\\\"\\\",2):f(\\\"\\\"{9\\\"\\\",2):f(\\\"\\\"}NKyb7bibhIR5?*ItPaubQ;sXO*bU1ye<k-t+1ye<4bpOQ;7?nDUIS4yb9.7\\\"\\\",2):f(\\\"\\\"{4VecU1VaoM+UN|:+*6ekae5tbVaoMab13eHbPaC\\\"\\\",2):f(\\\"\\\"}DzRM>z?uxz@\\\"\\\",2):f(\\\"\\\"{EPK\\\"\\\",2):f(\\\"\\\"}Z0rN7=@Hl|eGS2:+e5tuTa0b4b4q0.AaTny5mbebyzPaQae\\\"\\\",2):f(\\\"\\\"}xbVa+T67+b\\\"\\\",2):f(\\\"\\\"{bEaE1UacH,y4X,Xbrxz:oY>txCtTavD@-O+ShkIGgh9=@8bCtWaxr>aQaVsWLyw054b|bE^127^\\\"\\\",121"));
$write("%s",("):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^32^[2fha\\\"\\\",2):f(\\\"\\\"})3(f\\\"\\\",2):f(\\\"\\\"{#v3rga(f;)0,73-^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'ba6riOCEcZB3fN*,*,QaJp?Kvkws055g,bJn3bWabb21U5qZCY7b.vmueQ\\\"\\\",2):f(\\\"\\\"}p+w@LBoRa/qb\\\"\\\",2):f(\\\"\\\"}5x?9\\\"\\\",2):f(\\\"\\\"}QXKNwuhcow+A1HrdbcbTaM|NkJNSrAsqDcTP,xbNat*Mwa;fFa;Eah,K1PaAa?E<1xz0Lnv1qsVe4/b>;8blbPaoMgY7b4btb\\\"\\\",2):f(\\\"\\\"}usqlu\\\"\\\",2):f(\\\"\\\"{0.b6@3q\\\"\\\",2):f(\\\"\\\"{60su3a?ctufbvbShJOW>JdGsibaA|bW/9;.*;h+1\\\"\\\",2):f(\\\"\\\"}1VwNab\\\"\\\",2):f(\\\"\\\"}/bNab\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}1JCfbcz4j,bcb>kb\\\"\\\",2"));
$write("%s",("):f(\\\"\\\"{vbjP=jRaXa@?xbxs=oGT1pKH-005Vfy05Jjb1bFzxsvb.b679qo\\\"\\\",2):f(\\\"\\\"}vbebF0Xw.KC6H6TaSnc.k.HL4?*bibqYPpDa0bFaZ/TDQa/bQByb<aWrvbA1FaMAKC*2.bWrib?aSY<rp2L2j7v4\\\"\\\",2):f(\\\"\\\"}CRa82s+/p|:>ap2hbn/9q-sbqFD86e9cE3go+b5b|yPambxzhb7bU6E/@aI679vyz6bbY?HI2b0bw-5Uzb6vp3p.Bak|<t8x8bb8BHiAs|gbEG\\\"\\\",2):f(\\\"\\\"{rfvWaZavba2TambBpl\\\"\\\",2):f(\\\"\\\"{aSrl0Q\\\"\\\",2):f(\\\"\\\"{bEanwHTNnvbU3ZaXa*b|rVLXL6>\\\"\\\",2):f(\\\"\\\"{1>asM|VgANayb29Rsovc.=a*Tz<n\\\"\\\",2):f(\\\"\\\"{55:gd,D2fvLvH=87o;1T/9M+YKWKx0Ss1T57tbDp\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"}J+@R0Q1TSspt.i:Y9bDaO7b:a=a56\\\"\\\",2):f(\\\"\\\"{b|12|rXd6|bQabbY|8b;8q|vbjbT>s5n*o/DniR+bmbNsl,,be<B.nLcfb2FO:\\\"\\\",2):f(\\\"\\\"}B1xN64vUY*Q\\\"\\\",2):f(\\\"\\\"{z/9FZ-?BpDn>5g7XnFi>aDaQZabxXfbFa/X8J<ztx:PLp-hkZ6bOzEt?aUWbb@J.b5xMAYfT4gbeGczb-b|\\\"\\\",2):f(\\\"\\\"}Pv,kNr/\\"));
$write("%s",("\"\\\",2):f(\\\"\\\"}h*R45*Dvov6>eB1wOyOaYaAaF-1ulbL*Aa1T|N>yWaqOj5e|GMWa-bvy+9i;>1,o<,Raj61T\\\"\\\",2):f(\\\"\\\"{bx+UabZvo>a;VHN,*7s5N2.Ta@9^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'3ccakou3a<a/b6*M;n\\\"\\\",2):f(\\\"\\\"}t9x+ut7:5B910-xUbb*-5xAF+GA35Ni9i-x95N4b=a/b@SaNHfxdkb-?\\\"\\\",2):f(\\\"\\\"{y3ggVUaH-vs\\\"\\\",2):f(\\\"\\\"}b@oM;jbZ6>nH6TaGwiuf=D-PvSghbB;=aVvT\\\"\\\",2):f(\\\"\\\"{/.GGk4c*C,A|lbParNE.?z?*P|\\\"\\\",2):f(\\\"\\\"}07bQslK1*u+JpefHo/z|bgkl732.b6b2zuNg*WG:?.-rNX-4b1*27qWp=<a5bFa\\\"\\\",2):f(\\\"\\\"}QoOSnsVPDWrnL.4M<RaXvOtShJOcdNa,w,b>aYBYaGLCc|\\\"\\\",2):f(\\\"\\\"{Wa|1S/K88XH8A9fb4wRaQaz?.b\\\"\\\",2):f(\\\"\\\"}5+b6PQDUs"));
$write("%s",("GadR3xe8f<ATM\\\"\\\",2):f(\\\"\\\"{dzShAq5*Htzbr|kd.0RMA3+bMv:onr*qE\\\"\\\",2):f(\\\"\\\"}oO3bXFEs$6e5a.b>a-\\\"\\\",2):f(\\\"\\\"}wbeotv0b8ba11b-b2b<pU;bQm50b\\\"\\\",2):f(\\\"\\\"}q.b-bM|\\\"\\\",2):f(\\\"\\\"{bA9OzE3cka.b\\\"\\\",2):f(\\\"\\\"{rNga.|7q3e1c>az???;NqtGswb,bhbRavkjV+QdRq9246bw5s5GUU0\\\"\\\",2):f(\\\"\\\"}k,->AefgyFrQv3AAuwbT-tbA\\\"\\\",2):f(\\\"\\\"{QavbMrhp18u8bwn-I9yEd3@1FsfvFnJvAFWazbb\\\"\\\",2):f(\\\"\\\"{6bE8|\\\"\\\",2):f(\\\"\\\"}lb\\\"\\\",2):f(\\\"\\\"{r/b.bhr<\\\"\\\",2):f(\\\"\\\"{/bQT6bfW<\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"}?*2Eajzk.fWzdnpl6BKNkp=?U2burQa2bX0A\\\"\\\",2):f(\\\"\\\"{9+DS6yorgUIumq2r5*lb6-*q\\\"\\\",2):f(\\\"\\\"}DZsAqzbaR6b*5UaM<\\\"\\\",2):f(\\\"\\\"}?.6ega2b6bwPv4a+cXFebcbk.Pa|ub8a71bpSfW<\\\"\\\",2):f(\\\"\\\"{MAEauxQD|tzvX><G1bXMX\\\"\\\",2):f(\\\"\\\"{>ZgV*\\\"\\\",2):f(\\\"\\\"}ruAv2bfW<Gw-vfCs.ADw6bbQRvRaS,,vI<3bDoqZqUFaxb\\\"\\\",2):f(\\\"\\\"{b8vtv>,,v"));
$write("%s",("Prnt5vO?-uld1bbb/vYaib7tI9tbEa<aNaccHSAq??cT6g0v+A>|=t?abjAFWaiBv:gUAAXaYfS<D2@k0v+A?aRaXatb5SbC*b6bwEjHOH(ba7kIvZIvba7ZI.da,43?4[ha(f;)594A4.ia(ntnirpnt41da652t4.ba)T5[97[97[v3lGa\\\"\\\",2):f(\\\"\\\"}>tvAFWahb.\\\"\\\",2):f(\\\"\\\"{j4hr?LS,ld,*6b.vJvrKs?:*/b@aMvA|XaYfyb;1DAoOE\\\"\\\",2):f(\\\"\\\"}4U*5rC.v)>e+a7AcDBv|NX\\\"\\\",2):f(\\\"\\\"{o,mwUaM<.KFsrvpv3rBwLpf4Lpmxg3aCc.@w-wb6XO:md8BAoCc0b-YVa3b+,GaGSOaiMjk\\\"\\\",2):f(\\\"\\\"}uzbA?>zy\\\"\\\",2):f(\\\"\\\"}eb2b-u.bOavb1b9Wi3BC-uZMO5CajTm5qseb+b0p1sHY,b*5@53ioIR4V+bu,*cOShaO<5\\\"\\\",2):f(\\\"\\\"}u:5g675L//b15Py.5x\\\"\\\",2):f(\\\"\\\"}?-xb@CZBjb|blbHZy7Ya;Nx7fQXEjF|b-?X\\\"\\\",2):f(\\\"\\\"{l9X\\\"\\\",2):f(\\\"\\\"{EofbubEP:oeH\\\"\\\",2):f(\\\"\\\"{K2*X+GaGSVaupjWTizEi78bqgjkI6pBZ,Aan.+>C00HqU|6e2b8wEP:oO.JdnUg<tMxtN?,yJtn.3016K,7fx7mbj7y;eC8bBiQa:gO7>5-3Foc\\\"\\\",2):f(\\\"\\\"}"));
$write("%s",("Xa2C:P:o.ixu>r2tQaO+vDQank56ibqIywlt||.K+b=ao+ywTaf;ejSSKYtb*b@>WtS2tbZUaEb7|\\\"\\\",2):f(\\\"\\\"{b2bkx+bXLF39sB.Wa3bHVpoOa+FD@;N.Ktlx\\\"\\\",2):f(\\\"\\\"},*8shbQn.E:@S,e+lbJvX1Mt5bcTLZ1b6*I<QaQwnHAadXao>a216b,XDY2zib\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}gb=D>VQww0rqkbDrl9VrXnubLndwej2bebab9bQaW<wpw;4-Vfxa2bn;Mx\\\"\\\",2):f(\\\"\\\"{bqzs;ybTawqYCxbS$Y[v3aadhO:C:Taj4xbRa/sx+P:N:f;\\\"\\\",2):f(\\\"\\\"{;OrcQRv9bvg3b>Aybxb/ztbslvX79eE/sw+s;bu.KCE8/ybEyu5FZWa0-+D|;oi|UEax7n/o0CoqzU6d\\\"\\\",2):f(\\\"\\\"}b\\\"\\\",2):f(\\\"\\\"}|;xbEa4b4bWaYhab,bqgOa,yTaj4cvWat6u6vqj4aK8-H<zqv+0;8*qQ39EaybPa,yTaN;u5gG:or=F|Ea790|9bU6ybEyb;79I6k.xbj5w|Qa=CR+i8VaZaWH-4c.Uaf<3ve5s?NTYazXWsBiLz8s?pjYx>f+dby3F3Ngcb/wW>412pDan-dbTv-EHTtbSh\\\"\\\",2):f(\\\"\\\"{?nkRabQlt,tXzQ.3=i3cyOys=AxI.HDPaOn.bJ4wqv4jE=aup:=RaRaswcyGa5IWyWCzbPro?I<el"));
$write("%s",("jbYaygF7tbduRaQajLS,fbX\\\"\\\",2):f(\\\"\\\"{5b7+wbrpLAXaC,xGs?Rnd|Oadb;hrKUxCaXavr2\\\"\\\",2):f(\\\"\\\"{p=/x@Cj8q\\\"\\\",2):f(\\\"\\\"{ZazFQP5b,bWDF\\\"\\\",2):f(\\\"\\\"}1b1peb7u9<jY*Er:SQ\\\"\\\",2):f(\\\"\\\"}vhYG<K*8b?pDa8bitH6,6F-AaOay6Aaj3Va3bBa;vI6/b1UAaC3Ta;\\\"\\\",2):f(\\\"\\\"{Sas6C3nh/b=2Sa7bPa/b02ZaSG46eMaOaZyqwPCk1xLPFC;6/=aE8x=>aQa=V7Drj7DQ.jbits|**6bU6hb1rTa\\\"\\\",2):f(\\\"\\\"}.byAPRaE+vb<Okw64c.c96kb@ahkxZ:oMfDzAa*E<9pISMVat20bejf/7bQwY2-u.bc\\\"\\\",2):f(\\\"\\\"}VwibxbbqMviQ@agbf/c,6bntWHG\\\"\\\",2):f(\\\"\\\"},0>\\\"\\\",2):f(\\\"\\\"{Wy.\\\"\\\",2):f(\\\"\\\"}p,qQ/y+bDwu|b9bbw--bdb\\\"\\\",2):f(\\\"\\\"}.ubFaxE6rx=>aGU@>1Uf=jbDa+WUaybmt<aJH*b3b5b>aTzE\\\"\\\",2):f(\\\"\\\"{IXyB3.,Tg|N?=qgV5|91WaOrPq4oyBS1CalbT/1\\\"\\\",2):f(\\\"\\\"}bvpu>a0b<pSGVnEpGUi>Wf~bnurH1bXakbX\\\"\\\",2):f(\\\"\\\"{bYJ/?o8btbShKTWaE\\\"\\\",2):f(\\\"\\\"}:MZX*bhbXz=aib|bcjwvJ"));
$write("%s",("NWaDaYZwp9w,di|Oa*qm\\\"\\\",2):f(\\\"\\\"}>,+b\\\"\\\",2):f(\\\"\\\"{bAFjFD2kd,\\\"\\\",2):f(\\\"\\\"{.BS,KtAnwbOabbe1q44@:gJ4?P@wQ3aicnkbj8b@Jdb15kd.0mbwPV9XVrt;4fv?a;+mb2bQ;gShpqLvbDa**VN5v7uT*e5U@.QAnJ;QaFqPU@q<p6*vqH=:oR;>acO6-*qc>-bjpDa1b>a6-BaaxIvSrzb*D\\\"\\\",2):f(\\\"\\\"{.Xacl*bjq\\\"\\\",2):f(\\\"\\\"{bFnVN5v4b;/c\\\"\\\",2):f(\\\"\\\"{hbKv6b@ahx=v1bXajb\\\"\\\",2):f(\\\"\\\"{b>,2bdb5xBCDaQB86eOcEax9MpZR.Jmbi|z\\\"\\\",2):f(\\\"\\\"}sA+bjbdb94Ba4wpDVNRv<awbrqAsOyFa5:F+c8ShaOZ7EvP7ywTaAsH43K1KVa2.5oMOvb6vWLCt-@K/2brznwbbyrCa0RitQDg<Nayb?DZtMvLlsqmbs.*q<a1byDHpl|FFI>bo>x2|15t>2C=SWyMAo79yq4t,h9=@Ea+G=ARa9bBXEs,s*bnKlb6rs+eB\\\"\\\",2):f(\\\"\\\"}C=YY:zs4bVa+.:oE0t<@DDajDOaEtlu9bFa2|>amIeJdV:QZFaa;l90b<+j9cb.b5-SavbuhRa+P\\\"\\\",2):f(\\\"\\\"{Jq@QWi<kyRaU5zqCa@|As<a1wrDqArDVaZN0qS,7>gbShAPWLC\\\"\\\",2):f(\\\"\\\"}b\\\"\\\",2):f(\\\"\\\"}:"));
$write("%s",("hWaBK+b+wwsebNa4blbFal+Wygfe4\\\"\\\",2):f(\\\"\\\"{1o3MubBK\\\"\\\",2):f(\\\"\\\"}Z060*Qhbqw,b5\\\"\\\",2):f(\\\"\\\"}uw>YFa=onHNgnNo,sorL*qbAXnG>2VqMUMMOpuush-9x/w8B/wPyUMqM.EREjbtv-ba,4bEv,qeE3bebgo|blbubMOLqu=qqg2xTtUOa7LQwgoD\\\"\\\",2):f(\\\"\\\"}pr3b,r-E\\\"\\\",2):f(\\\"\\\"}4u=rKMO*:crSa6p@nvq3babrh=aqM7@<u.d,\\\"\\\",2):f(\\\"\\\"{=a+bXaeb=a+bWHzbMOIIqM2rF\\\"\\\",2):f(\\\"\\\"}>azbsz*6cea\\\"\\\",2):f(\\\"\\\"}NM<13anbQw.dHhtvTD\\\"\\\",2):f(\\\"\\\"},3>PsabJs2bW/CHZzmbf=go-UP7qQN\\\"\\\",2):f(\\\"\\\"{SaYhybQ-nLhbSatIUstIer;?fb?aBa.iOaZa@pBpnrI91Cc\\\"\\\",2):f(\\\"\\\"}y<qIl?ShKTe3g#aSa4q35H38b6B961\\\"\\\",2):f(\\\"\\\"{kvkbc\\\"\\\",2):f(\\\"\\\"{KKQaKYU;V6c0b.b5icu*9JC2|>aupz\\\"\\\",2):f(\\\"\\\"},v=aqv|tqJMv:\\\"\\\",2):f(\\\"\\\"{VQnpOaY*@,nNj2?Fpz*qG\\\"\\\",2):f(\\\"\\\"}P7wbO?:oLf0b\\\"\\\",2):f(\\\"\\\"}qLQoweo7QHsYf3bBa5b6bQwAD,bgy7r>FF=DaEa,Yv+kLsxxb+yP.qvi3UY\\\"\\\""));
$write("%s",(",2):f(\\\"\\\"{F3zy=eUtsovbNn4p5b>y5b|tqJBvNaybPtXaK,dXuNWa4vQ-ZaosaumxfWkpv0sA>yVaJleLOanHMfnN:o.rN<6bQwZaCAw-zb\\\"\\\",2):f(\\\"\\\"{\\\\\\\"\\\"),\\\\n(\\\\\\\"\\\"\\\"\\\",2):f(\\\"\\\"{ws,15b1u|NBvE0q\\\"\\\",2):f(\\\"\\\"{QD\\\"\\\",2):f(\\\"\\\"}b0B7bHpXK-|kv6bkb;z5b\\\"\\\",2):f(\\\"\\\"{rkb3XVfCak2eZhXxbuNCa9bZwL3Eu0*k3X*zb:*RaxbwpGs4Y;8dzhb32Pz+o3.kw;+MOSHp,2\\\"\\\",2):f(\\\"\\\"{XF=j5N@wEr8m9bB9DGm6I<4ygbcb<aeZdHArpO@Jq\\\"\\\",2):f(\\\"\\\"{zoJ1Y2QG@vhb|b7ba\\\"\\\",2):f(\\\"\\\"{6bF;uNmb-+/b|B|bFPZ,Y.T7\\\"\\\",2):f(\\\"\\\"{RPW8bDa0-ShHA=w5i7u8b\\\"\\\",2):f(\\\"\\\"{rJsHzhbNaNaZadq/b*/In5bm61-E8*oNgWyYVib<aib4bQqPCVa0-:oxzX1Z6tqUak*ZaEaWaoIkb.:7>4w7O<QL+:oxSibPauvytl9fW9qAatbX0bbSFFap,;\\\"\\\",2):f(\\\"\\\"{l+39qvUtzqjqR;Sho8LshX\\\"\\\",2):f(\\\"\\\"}9Z14|qoe|o5EacoHDFwgtm|K15|dTopt7m2Sh1G6bVquqF0DU?aJttulb4*GQkbxTz\\\"\\\",2):f(\\\"\\\"}dbiMQ,?EUa\\\"\\\",2):"));
$write("%s",("f(\\\"\\\"{TEt,b.JBD>VBKubL,UamuCAi/4JFaEsfbgbl71\\\"\\\",2):f(\\\"\\\"{l7Kt|<aRrj/y82mu937F*ReVcb79n3J@Jd777+dwh68/Fu3wh68bJVgbAwgNdbG8B\\\"\\\",2):f(\\\"\\\"}9udb8kuWab?wibGuPB9S**bQ6>X0eb\\\"\\\",2):f(\\\"\\\"}bAaj-s,r04jY*0:?aGaoW\\\"\\\",2):f(\\\"\\\"}uXHbWBa4*cPEaczF+-u.|Na;?*+fbkb.M.\\\"\\\",2):f(\\\"\\\"}:Q>5V9EaQsyrK1SKcz*06RSy<al-K-HVFVk3EaWzQa5bYa8bzGxGH>qIzxn,Qa,b3b\\\"\\\",2):f(\\\"\\\"{t0tMMIvCaVfK:5b9x=a-bhqt/npXa5b6\\\"\\\",2):f(\\\"\\\"{efi3\\\"\\\",2):f(\\\"\\\"}Cg<@Jnww**TX|8If\\\"\\\",2):f(\\\"\\\"{cb46hrtv\\\"\\\",2):f(\\\"\\\"}I7bvUMfw+M<nuDUBa+PpTlKFrv4VUNklKq2YfEUfhO|1b\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"{G*4sMT15C\\\"\\\",2):f(\\\"\\\"}gElbkqLfR.+bg4w02bp\\\"\\\",2):f(\\\"\\\"{b\\\"\\\",2):f(\\\"\\\"{;ve5vqINRE46\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"{EJQqvbsvd|xwP\\\"\\\",2):f(\\\"\\\"{j-|*@a*TgUSa@awblbCaJCtUrUpU8,@aZ/F9U5xbgbur0bDBfCvbQ/:z4JO.oA@yCabCX\\\"\\\",2"));
$write("%s",("):f(\\\"\\\"{g5RaUaCzAzMIxbab7?R.+v1\\\"\\\",2):f(\\\"\\\"{Oa2b,KcH\\\"\\\",2):f(\\\"\\\"{1@a5x\\\"\\\",2):f(\\\"\\\"{b*TMzXa0bCHc,22nwh-|<FP-@\\\"\\\",2):f(\\\"\\\"}v2k.ujFWqo+y-9bNICs,bAs:5/bNJptbqeoSF-bXaet8b2pxzvrBacoQ.-l|L*Jes|J+PqCbbg8\\\"\\\",2):f(\\\"\\\"{-rjdb=a\\\"\\\",2):f(\\\"\\\"}4Uzt+G.Qayb@RU9UxJv69<QPr,OY*,bV95ri3N60Ndb1*so\\\"\\\",2):f(\\\"\\\"}bpOShTQr*c.wbk1b11sjAA14vhbDyLG6=Ea*bYa2NhbGp\\\"\\\",2):f(\\\"\\\"}BmSAw7q3x-?6gC*fb8G@Ph4RM.q\\\"\\\",2):f(\\\"\\\"}b2beB4jhrZ0=j@y-b*btqCs1R5z8xEPBQ8rkb\\\"\\\",2):f(\\\"\\\"}s/y7b5Q94>agb?-ybVn\\\"\\\",2):f(\\\"\\\"{q<a>A-bO.pIg4x2=.2b.vNNk4NghrrL,btQ1v\\\"\\\",2):f(\\\"\\\"}o<uAoxqEqeC.@W0NrLrO+Aa6|\\\"\\\",2):f(\\\"\\\"{bybGp3Pkb1P|br|GaQ90lq>\\\"\\\",2):f(\\\"\\\"{L6HI5tBk>?arsQq@a7|k19q?,Jv;0bbZxxuhxibfb>xCp.-@*Shlwfb7uZavIVrEtkN0b98vbUGMzPaXaKJ5@QvTxCp4e0@kx5b3i<x|syy<anLSasg.+NI4b0Qg8Ua=C9bEqCNu*,i\\\"\\\""));
$write("%s",(",2):f(\\\"\\\"}bg<Xaur/b0sPvGaivmbfb/JqJ*bz*M\\\"\\\",2):f(\\\"\\\"{eb1=H1TavbRa\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"}:o*2hbWwHNX*\\\"\\\",2):f(\\\"\\\"{b5xab7bjbw\\\"\\\",2):f(\\\"\\\"}hbubYa*-6+8r0BYA8s:Pybw\\\"\\\",2):f(\\\"\\\"}9;>rDa29opI85\\\"\\\",2):f(\\\"\\\"}EGHDM|\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"},bOap\\\"\\\",2):f(\\\"\\\"{7IK1.b.bKC^127^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^32^[2fha\\\"\\\",2):f(\\\"\\\"})3(f\\\"\\\",2):f(\\\"\\\"{#v3rga(f;)0,73-c1Y:=\\\"\\\",2):f(\\\"\\\"{zoaIzbS\\\"\\\",2):f(\\\"\\\"{kbeLTaRaT<:\\\"\\\",2):f(\\\"\\\"}?2?M1yfK7I?*4a\\\"\\\",2):f(\\\"\\\"}Pdn,Nz<ShSt0-e2ebK\\\"\\\",2):f(\\\"\\\"}YCEoao\\\"\\\",2):f(\\\"\\\"}>2I9w|\\\"\\\",2):f(\\\"\\\"}ebb81zy6@a<96ONa1r@y;v2bBBMuzbrqeqybWa=twqT>0bx<o|S2r6CaUx98ub,:Lojbwb;\\\"\\\",2):f(\\\"\\\"}HsIN-ywb<N82mduN/bDr7olbuqkbYauNAav4dOR.vgzr=<|*Xa+bELIv=wPaqwkb.?Aaut\\\"\\\",2):f"));
$write("%s",("(\\\"\\\"{r,b3@@LlbjbNaP|qwnr7=eqZ0bqUnpxeBwbdb:oFacbqr>ajD3bA41uDv+CsALG2ElbCNejKC4bOawb|N1u6/\\\"\\\",2):f(\\\"\\\"{Klbf=ub.q.b9882Tx|b-@F3Pt7ta|Pa@adGbbvs9b=*Us|l*NYo*LQawb9sK\\\"\\\",2):f(\\\"\\\"}bb2*H|pN2bp3kbibubVLJ.lbUqi|Uahr=7/nfbfbQ|/1ebwqRamb1=2bOsYGzbYfxblb,b\\\"\\\",2):f(\\\"\\\"{tDa@DybU,.J7/EqA24b9bbbgbv:?MmvBadbd\\\"\\\",2):f(\\\"\\\"}Ral,3bOaM<D-Zzf>59c-\\\"\\\",2):f(\\\"\\\"}MCa07+bWav|E\\\"\\\",2):f(\\\"\\\"}bwOLu.zbzxBw\\\"\\\",2):f(\\\"\\\"{qBwD/x0+1vwfb0bk3Ba9-Eaub*1m\\\"\\\",2):f(\\\"\\\"{k2nuyz=apxF+DiS|QwUa*b1.zbWaYa*b=zwzdc4?,3Xn3b=jjb\\\"\\\",2):f(\\\"\\\"}b1b\\\"\\\",2):f(\\\"\\\"{>t6wbcbm0|bPjB7H.2C9b<a77L15b=>8s1rqJRa>sE+tuQ@JoDawbqDXilpR50lzJg:k:/DqBWEnwnuWyY:us:qhbnk5\\\"\\\",2):f(\\\"\\\"},b*b<p/pfb1bKo\\\"\\\",2):f(\\\"\\\"}bybPpwbnj|bmdM+zbw<dbtlnu2|VqSa77nk:*-bvb;qghwbnq*IBB=a0b-wv|1vybH>QpQaHzHIGq\\\"\\\",2):f(\\\"\\\"}4QwqD"));
$write("%s",("vpe<2B<pr3\\\"\\\",2):f(\\\"\\\"}bwbb8dw3bkbW57x|qvr7|;u0b5bMz4bLwJw1CU*7uubfb5>kbVaGa2>A7F|0JUISaFa94\\\"\\\",2):f(\\\"\\\"{d4p\\\"\\\",2):f(\\\"\\\"{dyb-bF9b6Tscb+r59CtJ4LtYa9bVaEae0h4,kx=8<4wA62b\\\"\\\",2):f(\\\"\\\"{bygrI\\\"\\\",2):f(\\\"\\\"{o2b:g,b9tA4OapDackbfbQt=abbKnIntbosBy/b6\\\"\\\",2):f(\\\"\\\"{Ou0DuBWuh:-l7H|ba.,bX\\\"\\\",2):f(\\\"\\\"{2rs5F4bulbb9O.4gy\\\"\\\",2):f(\\\"\\\"}*bUg2\\\"\\\",2):f(\\\"\\\"{<4Po8,c+a+\\\"\\\",2):f(\\\"\\\"}.B-nw8GdcjHpsWpU8,b?tX\\\"\\\",2):f(\\\"\\\"{9s\\\"\\\",2):f(\\\"\\\"}IY\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"}IYaBaWnu+cblbSaT,b3|\\\"\\\",2):f(\\\"\\\"{b6qsY-,q5r-w4jF3qt?a5pHByzOaSh>9,-@|\\\"\\\",2):f(\\\"\\\"{bns;>A>\\\"\\\",2):f(\\\"\\\"}bib39jH8wZacbb:l7Po?EszUavFdb*:Ea\\\"\\\",2):f(\\\"\\\"{bjbSa6+k3pB6bfI8/F0\\\"\\\",2):f(\\\"\\\"}kK:mEFue3E:dl2Bv|0bfbhCyuyBaub8W2xz5879I<H?eb:5S31b3e\\\"\\\",2):f(\\\"\\\"}:g-@<\\\"\\\",2):f(\\\"\\\"{b|<aoAab8irFvv+z>S>,\\\"\\\""));
$write("%s",(",2):f(\\\"\\\"{935H433FtbOa1vwpC,OnY*HvA2LE1b7w-s;h.ul\\\"\\\",2):f(\\\"\\\"{czq88wV\\\"\\\",2):f(\\\"\\\"{T\\\"\\\",2):f(\\\"\\\"{bH@a@C+bwbPaD\\\"\\\",2):f(\\\"\\\"}9bkbWaPjQa6*F9mbbvab<aGg>@ab<ztbDaCa1qjbno+bZB6bYzym4b7bcbO*y\\\"\\\",2):f(\\\"\\\"}55A?tb8bKfcby|*yJvdb7bhb6r:@n;NaEae2,/N6t@Ottbp?5s9;Sy0bUa5b46,6hpwy\\\"\\\",2):f(\\\"\\\"}bkC,r<a>kU1IuE0tsK,6b3gmBSsC0N*-|NgFa\\\"\\\",2):f(\\\"\\\"}9*bUa;>Z|W>kC.Eabs.=wc*5bvb=aDaRaBagb/9;ETpFa:\\\"\\\",2):f(\\\"\\\"{Zzqs7z:tX\\\"\\\",2):f(\\\"\\\"{j2rvZa\\\"\\\",2):f(\\\"\\\"{1lb8bxw;<o;p2/.Y.X7p>o@U7rBShM=C4ShD:<a51<a3blbc-n/abL2A3@A5b5bP=Y:??ZaEtymubXal-I+2bCsk+,q=BVal|?p2bybWv2bu7kbWyHwup/zXaWz+qh-Y>@tOa5.67|byhovYhr<vrbbUaD=H4YaY1x\\\"\\\",2):f(\\\"\\\"}KuHz;Dyh@|bC\\\"\\\",2):f(\\\"\\\"}bdB|7t<\\\"\\\",2):f(\\\"\\\"}b/./BbCRa,b7bGpEa6b5bTpY|6b+bo+71Gws\\\"\\\",2):f(\\\"\\\"}nuurKCB36b/\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\""));
$write("%s",("}bC6v9@a*\\\"\\\",2):f(\\\"\\\"}/xND?sQaeb?eY:OD9qQ0G\\\"\\\",2):f(\\\"\\\"}o|>a2kSaPB*95bZaYf6bK+7bfbEpuqab9zAaxBK\\\"\\\",2):f(\\\"\\\"}|z1bybVa.bsto0Cv1p.|+bCagbLz-lf:p@93n@93l>Wmrz/bUaLsWa.bq\\\"\\\",2):f(\\\"\\\"}2kWacb+9xbN7dByb@a3bFa=v/bZt\\\"\\\",2):f(\\\"\\\"{bt<ebD|X8iboqmqEv@ajkCaAa\\\"\\\",2):f(\\\"\\\"{bgbxbB3aj0C.C5-Y:Va>Bur:CZ?Favblbt<;,>yr0/w,bWag/hb8b|b?a|;Tafo?aVabCZ?n+<aablb-b-bBaao\\\"\\\",2):f(\\\"\\\"}BeC<acCwbP,I1:5NaI4wr5\\\"\\\",2):f(\\\"\\\"}VaFaU@NaM;D|n;p+vb3v0b@2x|cblydzwbAzFa<aU;RaPazbizCnBahp:\\\"\\\",2):f(\\\"\\\"{lbcb=aNaVpsqc.g,KA7\\\"\\\",2):f(\\\"\\\"}Xa5*+5\\\"\\\",2):f(\\\"\\\"{xQaRa<acblpy3lbA\\\"\\\",2):f(\\\"\\\"}Da\\\"\\\",2):f(\\\"\\\"{oLu<albe9rvQamqlb+bc,lbss>a1*\\\"\\\",2):f(\\\"\\\"}bgkY13bmbNajrdb.bOum>E5o>l<m@ab:olb2xtuSakwzb?asqFaN7>a*bTpeo*\\\"\\\",2):f(\\\"\\\"{.4Ba.bky*,AaDayhQqSaUjOrX\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"{bRaebo"));
$write("%s",("i96?a:uRa1=|tTaswzb>az*RawbP\\\"\\\",2):f(\\\"\\\"{*bJnz<i-?7Y-Qsg6eb65<af7i|+bi-/vCaF|DatwOy.0y3o|t>N|6sR.4bR+zbhvEp7biu\\\"\\\",2):f(\\\"\\\"{d<jh>3b=afbPa.uFv?a4b\\\"\\\",2):f(\\\"\\\"{bC|jkbqdznoQav|t|b@0bo-C|r3J?597pl3j3F>=ahbFuxbF\\\"\\\",2):f(\\\"\\\"}*q4jm6Oz77bzubV35bv+QwI;3bPaVa+bfhsx3b9-.bXaQ3M.P4WaY*7u8z.bvpcl|<ArFab\\\"\\\",2):f(\\\"\\\"}9333W7Y.n>j<ybOaA?\\\"\\\",2):f(\\\"\\\"{fwl|+E?nuz9b+wb?rTa7bEq7?1qi|btq|d>tz1?UaR+.4f\\\"\\\",2):f(\\\"\\\"{n8p3x*n+qqp,Iuabi,5vZahbTaO31bE9\\\"\\\",2):f(\\\"\\\"{bN<EaVa\\\"\\\",2):f(\\\"\\\"}bT9ettbc>kvzbVaOaabmbpzFa5oOao|dbxb?w=u5us>0bC>|bhbE.Vajbeb;;SaXq?2gbe1y+*b5/cz671/k+n\\\"\\\",2):f(\\\"\\\"}jbZawb\\\"\\\",2):f(\\\"\\\"{sGaI/\\\"\\\",2):f(\\\"\\\"{b0bhbN<x\\\"\\\",2):f(\\\"\\\"}|b.w9zb96z4zk3i35b283je3l7C9,b-8h*b-DaQaiu1boyZamb\\\"\\\",2):f(\\\"\\\"}bzyShu-ibX0\\\"\\\",2):f(\\\"\\\"{:;t9t7tf\\\"\\\",2):f(\\\"\\\"{-4Fax88bub"));
$write("%s",("Sx:8rt7bur<aYa-l83j:V7G5Y.m<d:c|o|zbnsubd,d|ibxg>\\\"\\\",2):f(\\\"\\\"}WaHzSnP/YwM\\\"\\\",2):f(\\\"\\\"{S2AaO=OaNartKx/b6bebp2*bgb2->aQq-blx*tRatwm2D<.rjpfhHti3VrZa-bR,Qxp2NkPa\\\"\\\",2):f(\\\"\\\"{sI<s\\\"\\\",2):f(\\\"\\\"}byp<h4S|6rr=|dI4Y|.bSnFuBa37+bNaI<*bPzPa>kuoFwBr@\\\"\\\",2):f(\\\"\\\"{ub\\\"\\\",2):f(\\\"\\\"}9db?ybq5vd1jqaoXqZz:o7\\\"\\\",2):f(\\\"\\\"{6+\\\"\\\",2):f(\\\"\\\"{blbtbu+Da075b.babz\\\"\\\",2):f(\\\"\\\"{wqNaNg1bnpU821Da-bwbZaj7u93bXz\\\"\\\",2):f(\\\"\\\"{b*w9b=al9<\\\"\\\",2):f(\\\"\\\"{>1bj-dTxJ.F4*8u*,bLl,dPqWa0b\\\"\\\",2):f(\\\"\\\"}u\\\"\\\",2):f(\\\"\\\"{bupu31bl8|rlbW|cb:ol7OuF5S7u\\\"\\\",2):f(\\\"\\\"{x\\\"\\\",2):f(\\\"\\\"{e:mbi/WaC,Saw1o\\\"\\\",2):f(\\\"\\\"}Pa>a5umuDayvcx>aSamdcbtb8zh4lbfbQr5bzb+brzDaNa57Et>axbyr-/jdgbQ66b-btu3bCcax*:Y*c|8b4yj4U1L24b8b@\\\"\\\",2):f(\\\"\\\"{qgiyf;\\\"\\\",2):f(\\\"\\\"{bvr*t4b4yG6B:hxQ2r4duyd4pYaSaRat6b2X0Rav+xz?a\\\"\\\","));
$write("%s",("2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"}J:b\\\"\\\",2):f(\\\"\\\"}=a\\\"\\\",2):f(\\\"\\\"{byzwbl4Sh=lhbJ*Y,Z,r5zq8b76L/X0Panyjjyw1555?9j2xz.hP/wbu/G6T,vyEtfbJpY1XaW89b140:Ea.:Ta-ydbl1>a,8Yafb\\\"\\\",2):f(\\\"\\\"}b3bv|8z<u*b7bQpS26bQacr-tQatlZ1Y.p1s1V\\\"\\\",2):f(\\\"\\\"}5393u123bbtbXa*\\\"\\\",2):f(\\\"\\\"{a3jblbab4b6bpoNwKq4\\\"\\\",2):f(\\\"\\\"{?nstc7prV387<xDa,bX8Faubb|*b-bOa|b:oQamb.bcxA.9b9sCaabwba6lb0bk*F+\\\"\\\",2):f(\\\"\\\"{b/v,b=aWaFa\\\"\\\",2):f(\\\"\\\"{b/\\\"\\\",2):f(\\\"\\\"{Xv2bP7\\\"\\\",2):f(\\\"\\\"{bj7dbRa\\\"\\\",2):f(\\\"\\\"{bw0sgJl\\\"\\\",2):f(\\\"\\\"{,8bzbEvtbu|swvb8b3oM4abFu8zBa;upoVpCadbb1kbBaTx4jgwr.uvK+5b:-h4npu,Etkb\\\"\\\",2):f(\\\"\\\"{,kb<anw<a/wP4j25sxu\\\"\\\",2):f(\\\"\\\"}wWaTa:oPo.wo*m*3xhpSaE\\\"\\\",2):f(\\\"\\\"}|b44S|1bmbV-pol7bbubmwg/WrAvJ7*b7uk\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}u*bZ+DaibA\\\"\\\",2):f(\\\"\\\"{xb1pW^127^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\""));
$write("%s",(",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^32^[2fha\\\"\\\",2):f(\\\"\\\"})3(f\\\"\\\",2):f(\\\"\\\"{#v3rga(f;)0,73-c1aWaLndb4y8b1xJd:o*\\\"\\\",2):f(\\\"\\\"}C,w\\\"\\\",2):f(\\\"\\\"{b/73w\\\"\\\",2):f(\\\"\\\"{q1t\\\"\\\",2):f(\\\"\\\"{H513h,tbSatbWa@aib6b6p>ai3Fa=7EpEaDaYaqzUsO.ibTsH|Y|Yw8bkb7bWa?aOazbi3fbU3s,j2c6/b>a9qzbx7QaCc4bmp16xb\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}=we+bzTwZz/qe0xbWwyb\\\"\\\",2):f(\\\"\\\"}bxbaojb=2mv<ac.t6/b=aj3ws+6Sact?,<sVaC|w6Wa\\\"\\\",2):f(\\\"\\\"{6xzq-Z,WaSalbKuj4vs=aX\\\"\\\",2):f(\\\"\\\"{hb6bvb:oR*o|I0Va:o2-lb+r7blbgoEqkb4p|6s|4/mb@a2|;hE3SaWaRaqwlbhqI*UaAaSae2SsSax2/bTal-Aa8zzbib5qp.YaQ37bBaPwI3gb0|>ocboi6p+b.i-v:oG-E-OaYww\\\"\\\",2):f(\\\"\\\"{IxD5Gxw\\\"\\\",2):f(\\\"\\\"{Exr1Cx?a+bk2\\\"\\\",2):f(\\\"\\\"}zYae18,VyXazbCpv|ub3b*ofv6rFaNai3co82@a*b?a7bfv\\\"\\\",2):f(\\\"\\\"{*8o9b\\\"\\\",2):f(\\\"\\\"{b5bb\\\"\\\",2):"));
$write("%s",("f(\\\"\\\"}|b7|Ya\\\"\\\",2):f(\\\"\\\"{brsQwhbfbtb6-q.|b|vcz+bnqRa1y1b/y-y+yAaTaLz\\\"\\\",2):f(\\\"\\\"{b6bRaNa9bgbUaS|po\\\"\\\",2):f(\\\"\\\"}bC0>w+b6bfb+v*b1x?uVaTx1b8wc|UjXaEaQaM+3b@2SyzpRaE\\\"\\\",2):f(\\\"\\\"}9bCa/vNwUacbu3G2E2C2VaA2?2=2;|Opk-0bK\\\"\\\",2):f(\\\"\\\"}A*EsRa?aVt6m/\\\"\\\",2):f(\\\"\\\"}vb>aOa.berOaxbvbTaPa@,Yf,\\\"\\\",2):f(\\\"\\\"}*o6v|bXa|b6b,|bjcz-belVaPp\\\"\\\",2):f(\\\"\\\"}0ubczp\\\"\\\",2):f(\\\"\\\"}/\\\"\\\",2):f(\\\"\\\"}bb.vUaEaqqSa>a7bKfZ\\\"\\\",2):f(\\\"\\\"{FnZ/0*ty4at1X.o1-lT\\\"\\\",2):f(\\\"\\\"}Y.3,a/XaV-B.Gz?aYahptum\\\"\\\",2):f(\\\"\\\"}Bt1t7bDa.\\\"\\\",2):f(\\\"\\\"}r\\\"\\\",2):f(\\\"\\\"}@w=a|\\\"\\\",2):f(\\\"\\\"{B|e\\\"\\\",2):f(\\\"\\\"{CyNaab8pd|8b+b@a-bbtF\\\"\\\",2):f(\\\"\\\"}8rtuubxbFan.z*2b9b1b/|EoQaFa8bEa/vgx0*>\\\"\\\",2):f(\\\"\\\"{jbL/\\\"\\\",2):f(\\\"\\\"}x;pIszb\\\"\\\",2):f(\\\"\\\"}b0pQadb+rcbkbAa,bDa*bUj2rh*Oatb?z.tcx?ajbAa\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\"));
$write("%s",("\"\\\"}\\\"\\\",2):f(\\\"\\\"{,<hv2HnH1RaZa+b:op\\\"\\\",2):f(\\\"\\\"{upkb;.vbYa6bib+bUn/bT|/\\\"\\\",2):f(\\\"\\\"}DaDz8bAa\\\"\\\",2):f(\\\"\\\"}bfbCaMxTaJ*/bVacbebAambYwnptbaxab/bV/UaT/G0E0Ea:oNa,b2bc18b>1ubCa2b1b1bF+Ba=jDaUa20>aTl\\\"\\\",2):f(\\\"\\\"{b*o+bZag1-bSmArfbhb>\\\"\\\",2):f(\\\"\\\"}Dab\\\"\\\",2):f(\\\"\\\"}tby0Fa-bP0\\\"\\\",2):f(\\\"\\\"{bYzI*Y.R\\\"\\\",2):f(\\\"\\\"}2,Xun14,6,W\\\"\\\",2):f(\\\"\\\"}OuucYa:ofxhb;0OaM05bc-=awbwqFasgubOaAw>aFzN0VfVa1.Qybbbbg0BaTlmbS/b0ub7babubi,y0xpZab\\\"\\\",2):f(\\\"\\\"}G-6+|bsq.0:gu+c,xp|*7bsxeoTp-xdbXaxbzxw\\\"\\\",2):f(\\\"\\\"}vb\\\"\\\",2):f(\\\"\\\"{.ZtScabgbwb4bv|2b.p3bTptc3bV/lb3o|\\\"\\\",2):f(\\\"\\\"}K+ubmb4bkqQaT/6-5s=jhbbbg-Eal|K/\\\"\\\",2):f(\\\"\\\"{bcb5-1bwbV\\\"\\\",2):f(\\\"\\\"{Mrgb>ambShjxmbCt.bEaPaKwt*D-8,ubibdbczjb:tAxAa8x6bTaXabz7pVt3x6-|oJ-mbGaYs3oqz9+6b1bebb|QqosSaPaY*Aa/bjbgbu\\\"\\\",2):f(\\\"\\\"}|\\\"\\\",2):"));
$write("%s",("f(\\\"\\\"}Kw*o.b>-eb5b+oShJxY\\\"\\\",2):f(\\\"\\\"}W.IbQ\\\"\\\",2):f(\\\"\\\"}ep5,5biblbYaQaPaFa|bz,Yamb8*1b?a\\\"\\\",2):f(\\\"\\\"}b,bFpub9\\\"\\\",2):f(\\\"\\\"{XaXa3b8bvbk-<aNryb?a@,5b6+Sm/bCsWa\\\"\\\",2):f(\\\"\\\"}bgbG\\\"\\\",2):f(\\\"\\\"}Ya:z9bxbPaZaPaab5br.hr1r=zec<aYnbbmbcbAa@aWa=aSa.bM*Tx<-.-AaZaFaebCydbi,jb*b2*/bEj4b;|V,=aSrRrS,\\\"\\\",2):f(\\\"\\\"}bP,eb?,=,=a.bSaab=al,q|Sy3gibCaQaeyabcb\\\"\\\",2):f(\\\"\\\"}bPai-EaRaNs2uAaPaWadc:o;heb*tdb/y7|Yntr1b.u7bLr4bNnKsibXa=azbOaM,4bNaubcbzb/bBafbbu1bUantVambl\\\"\\\",2):f(\\\"\\\"{C,2b+bkbQa9b@aEa2rBpfb|bvbSa=atb=ak|Cn0bdbn,XzjbUaYa=amb=aYa3eYaOu.l1,S\\\"\\\",2):f(\\\"\\\"}ZuX\\\"\\\",2):f(\\\"\\\"}P\\\"\\\",2):f(\\\"\\\"}gb1zy\\\"\\\",2):f(\\\"\\\"}*ytbybzbmbdl*btb.bfbopmp6v2bDa\\\"\\\",2):f(\\\"\\\"{b9zcb2b7bJn8b6buoQaBaEaNa|b@aUa=aXa:o=axb0b\\\"\\\",2):f(\\\"\\\"{booQaWaEacbTv1b@v6bDa@a|b9b+bT|abbbZaAajk0pwbUaM|"));
$write("%s",("@aN|,bib0bJtBiPaNa<w:wFw=a3b,*zblbp\\\"\\\",2):f(\\\"\\\"{ld>a3w0pSa.zWaUa8bOa*bVa4bg\\\"\\\",2):f(\\\"\\\"{u|YaYa<aOaeb/\\\"\\\",2):f(\\\"\\\"}-\\\"\\\",2):f(\\\"\\\"}M\\\"\\\",2):f(\\\"\\\"{*\\\"\\\",2):f(\\\"\\\"}OzqtYaDaubWaejAwgbbb-bCa,bPabb2bFi/bAaRacbubTaSambzb@a\\\"\\\",2):f(\\\"\\\"{*xqDzeb,bjb9sdb\\\"\\\",2):f(\\\"\\\"{*+b*b0*Ca*bTa**<a?aShd**b>aNaJykb<oZaDzzbZaUaPa1bwqOrnwct@aBa*b1b8b-wlbmb1\\\"\\\",2):f(\\\"\\\"}/bCatbc*kb=wbb4s0bVaDzwyfniiU\\\"\\\",2):f(\\\"\\\"}cp0lgiUuw\\\"\\\",2):f(\\\"\\\"{SuYuv\\\"\\\",2):f(\\\"\\\"{TzCvU|4y2bNzMrq|Sa0bzbwbNav|gbZa8x1brpsz6bbbwb-p6bLf<a8xlbnspuaw0b7b*bPaaw9bZa4bwbYaabab1bUx6b4b@aXa@aArbb3bwb5bfb8wu|\\\"\\\",2):f(\\\"\\\"}wGh|b8b=akbgbuf,bkbbbib3bZa8bSa/yybNa?aFa*b:p7sVv7pib6oQaxtTaUaibEadbbo?aRxSp0bjb9k\\\"\\\",2):f(\\\"\\\"}vNacbbbNaSa8bNatb?aCa3bcbqzBa2b\\\"\\\",2):f(\\\"\\\"}bbbabWa5btbgbFaOaWaub\\\"\\\",2):f(\\\"\\\"}b9x:o-d@"));
$write("%s",("aFabbYvcbVagbebtbebxbxb>ayb/bkbRaVaab@a4bdb-uvb+bPaebjytuMqZtLxqo@uYadwSqRrwb/brjhbcb/babXa8b5blbQa:owbFakbPaufjbPaUafbSaxbNgTabb4bfn4aRus\\\"\\\",2):f(\\\"\\\"{TuFxHxlbBa:oMvCa4b*bsqa\\\"\\\",2):f(\\\"\\\"{.pOzibTaDawt-bZadbhb>aebvb?aub|bYfIpBx2bvbbbebSa5beb1qcbFaybkbNa2i<a6b\\\"\\\",2):f(\\\"\\\"}bjb3b4q0b?a*bXaub8k|bWaBr2bQaTa|b4bhb>yxb<yYy0bAaab1vlbgbEaSxDpwbXaRa8bibbbKu9v:yEpcbYatbTyRyaqXaabkbswDa3b9yab7y5yAw?a6bNa@a.b:yhrCyAyRa0b0p4i:yjb;pAa6bsyhbYaZacv.bDa3iTa\\\"\\\",2):f(\\\"\\\"}uVaYaVa8b*wzxmb4jmbEambgbmbibBaWakblb5b1xZ\\\\\\\"\\\"),\\\\n(\\\\\\\"\\\"aQa\\\"\\\",2):f(\\\"\\\"}u@azb5o7bps8b\\\"\\\",2):f(\\\"\\\"{btbAa*bOambFv-b8b@apx-bSh4x2xix@afxejabQa=avbUaVa-u3bVa7b:oOuasDxbsOu,lYr,b6b,bct+q:o:tXaGuSaubgb\\\"\\\",2):f(\\\"\\\"}b6m:o8r-bab\\\"\\\",2):f(\\\"\\\"}b<aUa,bUaZaOa5bUa6vcb8bau2rYaXaCa8b7bTa*tNahx\\\"\\\",2):f(\\\"\\\""));
$write("%s",("}b6bjb:o\\\"\\\",2):f(\\\"\\\"}b<oPalbAa-bkbkb.dwbmb5b|bgb3b\\\"\\\",2):f(\\\"\\\"{bOaao0pabvbdb4bvbWa|bCaVtAaVa0bLqub2b8bwbibgbNaVa6pjb7b0bkbiucbgb5b\\\"\\\",2):f(\\\"\\\"{bzb7bbb7bgb*b|bab0bwb-uCa0smbjb1qFahbOa/b,kmbxbib>a:o|bAa;sebPteb.iEv0bSaebFabm<p5bNaXaoribwttbNaBaor\\\"\\\",2):f(\\\"\\\"{bUa?ayb.bmbabuvXaQakbSafbQa6b2vLsEa?a:ofv/bdbtu0bXa\\\"\\\",2):f(\\\"\\\"}b+bYabb6b\\\"\\\",2):f(\\\"\\\"{bubyb\\\"\\\",2):f(\\\"\\\"{bmb<u|bVa\\\"\\\",2):f(\\\"\\\"{tyt,bsr1b<p7b.bBa/b5b/b-bcb6bwbBaSh3s+bso\\\"\\\",2):f(\\\"\\\"{b3t\\\"\\\",2):f(\\\"\\\"{qAajbOubnVuQuYmdpcsOuhsdsfsgngsBbks\\\"\\\",2):f(\\\"\\\"{bAa|b*bbb1bfb,bSqVsTs*bEaCaPt0pebCpybgbkbmbts?aNn1rOaEatleb1bcbjbjkabib.bcb*bmb/b+bxb7bZaGt>acb0bluYacbabmjupyb3jRtjbybBa8b/bXa>aub7pdb*b=a:oSaUa|bkb:o9bvb,bRa7bNa.blbZajb@qYa3bFi\\\"\\\",2):f(\\\"\\\"}bqr2k3bTassOacbfbUasqqq3jRa5bDaybfb>a1bubNa\\\"\\\","));
$write("%s",("2):f(\\\"\\\"}bVatbfbTa2bjbEaUa4bwribWa4b:oyblbTagbZbdrWaNpFa\\\"\\\",2):f(\\\"\\\"}b@a;s5bwbCaShKrSq8b.bTaQaXaib:o3b/b:oYaeb.b=a4bPa*bFa/b\\\"\\\",2):f(\\\"\\\"}qbbxqybDaVawbwp8b^127^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^32^[2fha\\\"\\\",2):f(\\\"\\\"})3(f\\\"\\\",2):f(\\\"\\\"{#v3rga(f;)0,73-,#dbkp3bQa7bRaCa:o-bLqGaJq@a/bPa3b\\\"\\\",2):f(\\\"\\\"}bjovs+blbxb3jVaUaTaBacbmbmbXafbmb0b0bShyqXafngiapZrbpfpZofnfn;iToUaOa,bvbhrWa,bTaNa5b3b,b:oibQaYaFald,b4q4bubabdbzbkbzbMf>abq\\\"\\\",2):f(\\\"\\\"{rbc\\\"\\\",2):f(\\\"\\\"{b1bkb9b.rebzbNaprnr?aabVaCamdurTaYa-bWa8bFaSa|bdblbkpubQa\\\"\\\",2):f(\\\"\\\"{b.bUaSaVaubjbcb9bzbjbRazb2bVa2bfb6b?a2b>a+b5qwbub8bfb-b3bUaSh9oVaBa3b7b2b*q|qzq*b.bhbUavb@aIpvbvb\\\"\\\",2):f(\\\"\\\"}bbqsqdbkb\\\"\\\",2):f(\\\"\\\"}bKotb4b>a9b7bdb0bPa,babxb:o,blbUaQa>aib,bebVa"));
$write("%s",("rp8b0bWaBaFa+bSaEaAaUaxb\\\"\\\",2):f(\\\"\\\"}bebmb3bQo1p/pzb=a+phb*bBambPa0bEajbFaPaCambFa>aTafbibOaCajbhblbibkbcbibjbhp7btbbb|b2bLo|bmbBaDakb=a,byb|bSaZaPo4bQo.bAa0bZaDajbjb9bOaPaxb9b5bOa\\\"\\\",2):f(\\\"\\\"}bcbwbiiVoWo|lUo|lXoeniiinjniihnfnebDaFaDaTnebLfkbdb+bOaFaCawb*bCa<a|bZa:ogbvbNa1bGayo7b<a>adb/bSaXaFagb,o-o+o\\\"\\\",2):f(\\\"\\\"}o/bYagb7bAaFaShqbjbtcUagbYawb+dXabbQa<aTa\\\"\\\",2):f(\\\"\\\"{bwbEaeoVaRa>aFankzbdb-b3jeblbzb,bNa7bvbCaEahb<aCabb*bWgQaub*bWaQagbSa,bEa7b6bAaEaHl0nun:mkmimnnEf=mqm*n;aPmrm?apmPm<m:lznBmUg9lMmwbicPm;lhmqnEaSl=mjm9lwmemcmfn0l0lZm4acn9agian|lXm+lii/l/b\\\"\\\",2):f(\\\"\\\"{f-a|hub.h8a4mAmxmFm8l9aEaOa=m;m,m8f:a-b=m=aAa-a-m\\\"\\\",2):f(\\\"\\\"{mCaSlWlvm@a<a-b|e0mzmKlgmVlMlKlIlnmym:aCa|esm>aAahmRlMl9a6lNlAaVgDl|efmslHlUlBa-aJlClAl*bvbtb/b-a+bId<lOl=lFl@aDlHlSe|eBlG"));
$write("%s",("l?aAa9l\\\"\\\",2):f(\\\"\\\"{b7l>l<lFa:l8l6lHa4l9a|e5lxb8a+e-a1bLf8aEfpl8arb|eidfi-l-l\\\"\\\",2):f(\\\"\\\"}l3a:igi\\\"\\\",2):f(\\\"\\\"{l-fhiil<h7f6b-a+czbxbubHaqb6aqb3i4i2i5aqb-g-aff1bzb.b6fnbxbkiShHgFghgHfkhxhbkxjZj?a=a:i;d\\\"\\\",2):f(\\\"\\\"}h2kyiIjdh.ktcBa3a=h6g2iwb=fTjakFjBa?a9i6e|hrbLj?aJjSjviGjDa?aDj2b3b5iBf+c:g-a8f-b1jCa3aKa\\\"\\\",2):f(\\\"\\\"{b;atgwbccIa3b1bnj,b|b0adhyhdhzjRjvjCa9i.bbi?a?iyj=i;i@a9iyb3bBjyh2h>iwhwjBa>a9iPcsihghgsbubwbSh-a2j0j:a;b-j1b0b-b3aAa3a7b-aSh.a:b:b,byhlhxiPaUh<i@a3a|hwb+b-aPcbj/b8b1bPcxb;aBf-b;gZaWf|b.b5b-aTi,i3bDfvb|b6g5iWfMf3bgf;a<b:b3b-a8b6g,bxb2b2btb;ayhEhwiEh3a>a3a5anb-a3i/b3b4b.bHa8byb2bsgtbDfxb5b+bGgyhwhThGhlh?g8f6fHaoioiFaGaRh|fld4aogei/ach4a-aMfKfMaFa=aEh-bGh2h1hGa+bJd?h9a/b5a|fCcyg-bPaBaob2h6aKaMa9aMaIa5axb3b.b4b0bxb*htbLfyhRfwhGaMb5g2bzb;azb"));
$write("%s",("-b7fccJaWg?achlhCdYaOaVafbVaibNa=adhdh?a;aAgVaNaUaogchRfvbpbEa*c7b?a>aCaCa>anbJdubSczb=fIc?gyfwfuf2bsfNd3bHa?e-a-fGf:aIa+ctb,b:avbldub4bcb-btggcqgHaebdbJaGagfef8a1bxbwbtbxbUaac|b3bKffb/aRfggtbxc?f?a1aRf-a6a5bOf>azd:a,cNaOfwb.b;b>aHfob,c:a-a.b\\\"\\\",2):f(\\\"\\\"{bvbxb5a1aob,fCe2b-a:b1dtbHa6a/c2b/a:f-f;d+c1b/b3dMd-aDdBd@dmf/aob5a.d,d*d-b4b7eSc;axb+b.bbcZb0cbfJasdHa/aed+e0cGb/d,btb-b4aWbudpcgdLc=chchd6areOapc0cNb/a;bje/eGaHb5dedOb.a8aNd8aLdLa=a>aIaOaJapb6a+e5azb+cdcfbhc;aOaFdYd6aHaCa@aIaQd8aHa=a.cIbCbMd\\\"\\\",2):f(\\\"\\\"{cycvcocRapcXbocTa;b;bpbgbYdJaGbRanbQaJagbnbcb>dqc5dpbebnbOa8a0c4aJaTa5a+btb5bxbJaQa,c*cRa5a1bzc6aedMa0c3bldjd;aeded8ard5a6a5aedxb/btbvb2bxb,c1b4b3bxb1b0cocPa8aNapcMagdUc3b|b+b/b2b4arcFbnc4a=a?axbtc4aSbJcPbKckcic+bZb3b-bzcXbqcFb5aMa/ancvc+b+b|byb4a9cV"));
$write("%s",("bNa5aRb7cFbnbFbMapb2c.aMaFb.a4a5aJaOa-a-b|b-aeb5aicybHa<b/akc>a>aXb6aOb/a8a6a/apb4a1b.b3bvb4b1b3b2b-b.bvb4anb/aJaPa5a8a4a6apbEb5a5aBb,b9a4apbpbnb8anb4aGa=a:bJacb!5R1ca616R.ba~[2xha=s,y=z,54[54%.4[e6&yay,]99999[gnirtS wen=][c n3aea\\\"\\\",2):f(\\\"\\\"{)v]y3b&a(niam diov citats cilbup\\\"\\\",2):f(\\\"\\\"{RQ ssalc~5[~5qfa cdlnl3c/a;maertStnirP/oi/avajL tuo/metsyS/gnal/avajq5bdateg@3doa2 kcats timil.v3dga]; V);U5aC3ecaL[f6aa6hha dohtem?3e;4nga repus&3ecaRQ@3cgassalc.@6[@6ioa(=:s;0=:c=:i;)$5ajaerudecorp34[34eqa(tnirp.biL.oken\\\"\\\",2):f(\\\"\\\"{24bianoitcnufc:[83\\\"\\\",2):f(\\\"\\\"{martStup=niam^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\""));
$write("%s",("\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'>3(ba7U3vJ4vba7I4.da,43?4[fa(f;)5/6/#6[#6[#6[#6moa(etirw.z;)tuo.-@aba(q?b~auptuOPIZG.piz.litu.avaj wen=z|5[a7[a7;ca34A4.l41ba0j4[w5ada283m4[x5[j4fea1982m4.batv9[V:[?4:da12927[=8[V:[x5[x5vca04V:/5aR0Z0Z/512152353/2/2166263=4/3141726??:1518191:1/I9[.;[?4:da063.G/r9[/;[x5[j4Fda66957/da*6 .C[Z:[?4;da348Z:[A8[Z:[x5[57wca8457/ea1312aC[a;[?4<da423VF/C8[a;[x5[j4Fda200a;/YB[W:[YJ<ba1OV0>8[W:[x5[YJGca15XB/fa41310\\\"\\\",2):f(\\\"\\\"{9[[:[.[;ca92B8[B8[[:[x5[x5wv5/qa;t:\\\"\\\",2):f(\\\"\\\"}%%%%\\\"\\\",2):f(\\\"\\\"}fi\\\"\\\",2):f(\\\"\\\"}*-84OH2ca7786[86[Q8[x5[QPwba9R@/(a]i[\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"}+17\\\"\\\",2):f(\\\"\\\"{<84.;i:-i602\\\"\\\",2):f(\\\"\\\"{;i:911\\\"\\\",2):f(\\\"\\\"{;j:6323?[tA[?4:da550d9/xa(tnirP.tmf\\\"\\\",2):f(\\\"\\\"{)(niam cnuf;V4[;6[;6;ba93;[><[j4gca69mO"));
$write("%s",("/datmfY6[>8[5R;ca5847[?8[V:gca02?80saropmi;niam egakcapo7[O8[?4;L[1ga(tnirp[A[+6[?4;ca36(I/|<[j47da444l4.ba-W6[<8[i<[A?njanirp tesnw41ca21T9/la1 etalpmet.f6[F7[)L<l;/ga(ntnir|D[*6[?4;ca93SG/baf)6[)6[?4?ca11EG0$a,s(llAetirW;)(resUtxeTtuptuO=:sc5[C6[?4;8=/#BaC4[(6[(6[v3kdaS C&6[&6[*D<3=/ca&(?4[$6[G9[v3kba r=[)6[)6[r=[&6[r=[83)iaRQ margoP9[-6[-6[P9phaD : ; RW9[-6[-6[v3mba^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'>4[#6[#6[#6[#6[#6[#6\\\"\\\",2):f(\\\"\\\"}i=[$6[$6[v3lqa. EPYT B C : ; A36[36[36[y=[#6[#6[#6[#6[?4[#63ka)*,*(ETIRWs=[.6[.6[G@nhaA B : ;,6[,6[,6[v3lba [2cF4[+6[+6[T9oia: ^1^\\\"\\"));
$write("%s",("\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"' ohceI4[.6[?4[73kpastup\\\"\\\",2):f(\\\"\\\"{)(niam tniL4[164ca01?4[?43ea%%%%@4[%6[?4[%6[%6[?4[73\\\"\\\",2):f(\\\"\\\"}paparwyyon noitpo26[M45<4[<4[<4[<4[jD@hanftnirpD4[fa(f;)3D4/kaetirwf:oinu41ba2u4.ja>-)_(niamt4[Q8[<4fWP0gacnirp(C4-ia(stup.OIK4/rKajaM diov\\\"\\\",2):f(\\\"\\\"};)B3(ca11g62oatnirP)--n;n;)sn3a<a(rof\\\"\\\",2):f(\\\"\\\"{)n tni,s tsnoc gnirtS(f diov\\\"\\\",2):f(\\\"\\\"{noitacilppA:RQ ssalc[k4rga@(tnir>MblaM dohtem06x*3cl;abNcuadiov;oidts.dts tropmtNnra1(f\\\"\\\",2):f(\\\"\\\"{#(rtStup=niam&3kkaenil-etirwb8dva(,^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\"));
$write("%s",("\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'s%^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'(gol.elosnoc;)^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'73g\\\"\\\",2):f(\\\"\\\"}a^129^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\""));
$write("%s",("^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"' nioj.)1+n(yarrA>-)n(=fI3cva^31^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",2):f(\\\"\\\"}54,1\\\"\\\",2):f(\\\"\\\"{.^127^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"# qes-er(K7c.4cba^31^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"p3lg3fw3hla1% ecalper.j4dea^128^gXc/arts(# pam(]YALPSID^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^127^\\\"\\\",121):f(\\\"\\"));
$write("%s",("\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\".NOISIVID ERUDECORPA3cma.RQ .DI-MARGv3g53d|bNOITACIFITNEDI^127^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"[tac-yzal(s[qesod(^63^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"))System.Console.Write($^63^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"Put caffeine \\\"\\\",2):f(\\\"\\\"{(int)c\\\"\\\",2):f(\\\"\\\"} into the mixing bowl.^64^n^63^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");M3pva^63^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"Liquify contents ofE3oeaPour^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9)"));
$write("%s",(":f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'3w^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'4e\\\"\\\",2):f(\\\"\\\"{abaking dish.^64^n^64^nServes 164cma\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}^31^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");\\\"\\\",2):f(\\\"\\\"}/****/e3a^15^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"),s[999999],*q=s;int main()\\\"\\\",2):f(\\\"\\\"{int n,m;for(;*p;)\\\"\\\",2):f(\\\"\\\"{n=(*"));
$write("%s",("p-5)%92+(p[1]-\\\\\\\"\\\"),\\\\n(\\\\\\\"\\\"5)%92*87;p+=2;if(n>3999)for(m=(*p++-5)%92+6;m--;q++)*q=q[4000-n];else for(;n--;)*q++=*p++;\\\"\\\",2):f(\\\"\\\"}puts(s);return 0;\\\"\\\",2):f(\\\"\\\"}^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"))\\\"\\\",2):f(\\\"\\\"{s+=^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"00g,^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";for(m=1;m<256;m*=2)s+=^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"00g,4,:^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"+(c/m%2>0?^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"4+^7^\\\"\\\",121):f"));
$write("%s",("(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\":^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")+^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\",^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";f(s);s=^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"4,:,^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";\\\"\\\",2):f(\\\"\\\"}f(s+s);for(c:Base64.getDecoder().decode(^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"kaAREREX/I0ALn3n5ef"));
$write("%s",("6l/Pz8+fnz58/BOf5/7/hEX/OZzM5mCX/OczmZzBPn5+X/OczMznBL/nM5mZzBPu++fPPOc5zngnnOZzOZgnBMGAW7A==^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"))\\\"\\\",2):f(\\\"\\\"{c=c<0?256+c:c;for(i=0;i++<3;c/=8)f(c%8);f(^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"8*+8*+,^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");\\\"\\\",2):f(\\\"\\\"}f(^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"@^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");^1^\\\"\\\",4):f(\\\"\\\"'|sed -e^1^\\\"\\\",4):f(\\\"\\\"'s/^16^/^32^/g^1^\\\"\\\",4):f(\\\"\\\"' -e^1^\\\"\\\",4):f(\\\"\\\"'s/^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\"));
$write("%s",("\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"/^16^q/g^1^\\\"\\\",4):f(\\\"\\\"' -e^1^\\\"\\\",4):f(\\\"\\\"'s/.*/print ^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^8^nquit/^1^\\\"\\\",4):f(\\\"\\\"'^3^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")\\\"\\\",2):f(\\\"\\\"}^1^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")\\\"\\\",4):f(\\\"\\\"');\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\").split(\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",128):f(\\\"\\\"^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")"));
$write("%s",(";for(int i=1;i<a.length;a[0]+=a[i+1],i+=2)\\\"\\\",2):f(\\\"\\\"{a[0]+=\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",185):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\".repeat(Integer.parseInt(a[i]));\\\"\\\",2):f(\\\"\\\"}System.out.print(a[0]);\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");\\\"\\\",2):f(\\\"\\\"}\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";FORiTO UPBtDO INTn:=ABSt[i];print(REPR(50+n%64)+c+REPR(50+n%8MOD8)+c+REPR(50+nMOD8)+b+\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"J\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"+a)OD\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"while(!="));
$write("%s",("(S:length)0)\\\"\\\",2):f(\\\"\\\"{\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans c(S:read)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"D(c:to-integer)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 35 39\\\"\\\",2):f(\\\"\\\"}\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 24 149\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"interp:library\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"afnix-sio\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans o(afnix:sio:OutputTerm)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"o:write B\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");end;"));
$write("%s",("\\\"\\\",1):f(\\\"\\\"\\\\\\\"\\\")\\\"\\\",1):f(\\\"\\\"nsys.exit 0'}\\\\\\\"\\\")\\\"\\\",0)]]></xsl:template></xsl:stylesheet>\\\":s=\\\"   \\\":For i=0To 7:s &=Chr(32-(Asc(c)>>7-i And 1)*23):Next:System.Console.Write(s &n &Chr(9)&n &\\\"  \\\"):Next:System.Console.Write(n &n &n):End Sub:End Module\")\nput=s\nprint\nqa!"));
end endmodule