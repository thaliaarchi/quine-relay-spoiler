module QR;initial begin $write("%s",("let s=(\"Module QR:Sub Main():Dim c,n,s As Object=System.Console.OpenStandardOutput(),t()As Short={26,34,85,127,144,153,196}:For Each c in\\\"BasmCBBBCRE`F<<<<C<`C<B`BBD#CXwasi_snapshot_preview1Jfd_writeBBEEDCDGECB@IUDHmemoryDBH_startBDL|DRBAC BAJlACA4RB9MiCD<AERCA>D!BE@ABRCABRCABRCAJ!CE@ B-BB CACk:CvACqRC COBMADRCACRCADRCABRCABRC BACj:B-BBOBMADRCADRCADRCAFRCMM}CBABM~(BBBCBBB,BBBDBBB0BBBDBBB4BBB=BBB?BBB;BBB ...\\\\t..\\\\n..(module(import:wasi_snapshot_preview1::fd_write:(func(param i32 i32 i32 i32)(result i32)))(memory(export:memory:)(data :\\\\08\\\\00\\\\00\\\\00$:))(func(export:_start:)i32.const 1 i32.const 0 i32.const 1 i32.const 0 call 0 drop))\\\":c=Asc(c):If c=36:For c=0To 11:s.WriteByte(If(c Mod 3,Asc(614003.ToString(\\\"x8\\\")(1Xor 7-c*2\\\\3)),92)):Next:Else:n=(c>12"));
$write("%s",("4)*(8*c-39664):Do While n>127:s.WriteByte(128+(127And n)):n\\\\=128:Loop:s.WriteByte(If(c<125,If((c-1)\\\\7-8,c+66*(c>65And c<91),t(c-57)),n)):End If:Next:For Each c in\\\"<?xml version='1.0'?><?xml-stylesheet type='text/xsl'href='QR.xslt'?><xsl:stylesheet version='1.0' xmlns:xsl='http://www.w3.org/1999/XSL/Transform'><xsl:output method='text'/><xsl:template match='/'><![CDATA[sub f(s$,n)print(s$);:for i=1to n print(\\\"\\\"\\\\\\\\\\\"\\\");:next:end sub:f(\\\"\\\"write,format=\\\\\\\"\\\"%s%s%s%s\\\\\\\"\\\",\\\\n(\\\\\\\"\\\"\\\"\\\",2):f(\\\"\\\"write{-}{txt}{echo -E $'(\\\"\\\",1):f(\\\"\\\"\\\\\\\"\\\"with Ada.Text_Io;procedure qr is begin Ada.Text_Io.Put(\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans B(Buffer)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans O(n)\\\"\\\",2):f(\\\"\\\"{\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Chara"));
$write("%s",("cter\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"B:add(Byte(+ 128 n))\\\"\\\",2):f(\\\"\\\"}\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans f(v n)\\\"\\\",2):f(\\\"\\\"{\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"O(+(/ n 64)107)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"O(n:mod 64)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"O v\\\"\\\",2):f(\\\"\\\"}\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans D(n)\\\"\\\",2):f(\\\"\\\"{if(< n 4)\\\"\\\",2):f(\\\"\\\"{f(+(* 6 n)9)48\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{if(n:odd-p)\\\"\\\",2):f(\\\"\\\"{D(- n 3)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 27 48\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f("));
$write("%s",("\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 36 11\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{D(/ n 2)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 21 48\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 48 20\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans S(Buffer\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"STRINGz:=REPR226+REPR153,a:=z+REPR166,b:=a+\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"2\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"+z+REPR160,c:=b+\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"8\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"+z+REPR165,t:=\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"class QR\\\"\\\",2):f(\\\"\\\"{public static void main(String[]a)\\\"\\\",2):f(\\\"\\\"{a=("));
$write("%s",("\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"write(\\\"\\\",4):f(\\\"\\\"'implement main0()=print(^1^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"BEGIN\\\"\\\",2):f(\\\"\\\"{print(^3^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"echo ^1^\\\"\\\",4):f(\\\"\\\"'f(s)\\\"\\\",2):f(\\\"\\\"{System.out.print(s);\\\"\\\",2):f(\\\"\\\"}s=^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"389**6+44*6+00p45*,^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";for(c:(^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"#include<stdio.h>^8^nchar*p=(^15^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25"));
$write("%s",("):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"Ra#include<iostream>^16^nint main()\\\"\\\",2):f(\\\"\\\"{std::cout<<(^31^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"class Program\\\"\\\",2):f(\\\"\\\"{public static void M83abbSystem.Console.Write(^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"Quine Relay Coffee.^64^n^64^nIngredients.^64^n^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");for(int i=9;i++<126;)[3pva$^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",2):f(\\\"\\\"{i\\\"\\\",2):f(\\\"\\\"} g caffeine \\\"\\\",2):f(\\\"\\\"{i\\\"\\\",2):f(\\\"\\\"}I3b54rja^64^nMethodv4f#aeach(char c in(^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\"));
$write("%s",("\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")))^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^32^[2al3dp3c[2cs3c,3l[2k@3kqa^31^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")s rts(ecalper.h3eja^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"     53c4a SUTATS(egassem^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"rts(nltnirp(])]^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\".NUR POTSu4cba.C3dh3dX3bba[65bX4df5lga\\\"\\\",2):f(\\\"\\\"};)06xm3f$3loa)1(f\\\"\\\",2):f(\\\"\\\"{#qp]^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\"));
$write("%s",("\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'[p]#3sv3r23)ga3(f\\\"\\\",2):f(\\\"\\\"{#.33)ba7g4-ba5R4w23F&7d33&q7u53sda,4353.ma^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"' D ; EYB RCL4/v4+ja13(f\\\"\\\",2):f(\\\"\\\"{#DNEm4[m4ada. A~5[p"));
$write("%s",("4deaPOTSn4[#5e~5[o4boaRQ margorp dnex4[x4abaS*5[m4c2<[ba9i4[i4dba&#6[k4agaS POOL&<[77dba^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'j4[j4[j4gda&,)(6[<>cga. TNUO<7[s4bfa(rahcf:[(5dgaB OD 0?>[t4cca&,+<[ha9(f\\\"\\\",2):f(\\\"\\\"{#)A26[9=d4=[,6cqaEUNITNOC      01z4[a9c,5[U8dJ7[WFeeaRC .p4[p4aka,1=I 01 ODt4[OKecaPUq4[*I[5<gva;TIUQ;)s(maertSesolC;dYe$4Rra322(f\\\"\\\",2):f(\\\"\\\"{#tiuqn\\\"\\\",2):f(\\\"\\\"})652=5[qa^32^\\\"\\\",2):f(\\\"\\\"})974(f\\\"\\\",2):f(\\\"\\\"{#n\\\"\\\",2):f(\\\"\\\"})215iY3b8,ya99(f\\\"\\\",2):f(\\\"\\\"{#etalpmetdne.n\\\"\\\",2):f(\\\"\\\"})4208[.zX3ca02-Y[v3bda116~K[-L[j4ldamif+6[ga)30341\\\"\\\",2):f(\\\"\\\"}5[,6[j4l"));
$write("%s",("bat(6[(6c%a315133A71/129@31916G21661421553/04[04c(a%%%%\\\"\\\",2):f(\\\"\\\"}*+1%%%%811 -\\\"\\\",2):f(\\\"\\\"})48361(f\\\"\\\",2):f(\\\"\\\"{#j:+1 j@34[34cbawm4[m4cl4[l4cbaWm4[m4cba\\\"\\\",2):f(\\\"\\\"{m4[m4cva)(esolc.z;)][etyb sa)t=[#>[j4[~Jjca69m4[x5[j4lba,l4[w5[j4hla!\\\"\\\",2):f(\\\"\\\"})23(f\\\"\\\",2):f(\\\"\\\"{#~~v4[%5[j4hea(rt.o4[z5[j4hba)A7dda\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"};l3efa~~dneo3hra~~~~PUEVIGESAELPnr3ala~~1,TUODAERw3a63j$a(etirw;\\\"\\\",2):f(\\\"\\\"};u=:c;))652%%%%)u-c((||13jda#-<q3jda||i)3mhaBUS1,ODs4qka)3/4%%%%i(N4cx5kU4xPa2=:/t;2%%%%t+2*u=:u\\\"\\\",2):f(\\\"\\\"{od7 ot0 yreve;i-=:u;1=:+i\\\"\\\",2):f(\\\"\\\"{od))1(evom(dro=:t elihw?s;)s*45oi5vv3jd7dladohtem dne.s3dganrutern3d~aV);gnirtS/gnal/avajL(nltnirp/+Za|atnirP/oi/avaj lautrivekovniJ3d.4j[2cib\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\""));
$write("%s",(",2):f(\\\"\\\"};0=q;)]q[c=z(tnirp.tuo.metsyS;)0(tArahc.y+z=]++n[c;y:]q[c?n<q=y\\\"\\\",2):f(\\\"\\\"{)0>2%%%%++i(fi;48%%%%)31-)i>3c&as(+87*q=q\\\"\\\",2):f(\\\"\\\"{);87912<i;(rof;n)rahc(+K4r[2k*3&oa=]n[c);621<n++r4aqa0=q,0=n,0=i tni;N3&mc6axi4asdRbQeglxfvfZkRf<bedPd-j\\\"\\\",2):f(\\\"\\\"}b;agb-a|dzdxdRfGb8aqeRdYd5a\\\"\\\",2):f(\\\"\\\"{b2bFi;agb-epb>aqeRdHa>aJaRaAdteFbaeIfOa5aac2gO36f9aXG4aLa7a;a4a<aOhgmkdxd;aNa?c6a|eebHaFaIaebzeJaeb9a/a6a2dQbUe-f2a-f9aXG5d6cRbC3gQc-f/aof0fRfmh8kEf.b2e6aRa;dX-ogO\\\"\\\",2):f(\\\"\\\"{Fh;aTapc4aLcEexiof6amc<byg-f>lsbvh;CWfybxcxc>aGaUeAa2a6a\\\"\\\",2):f(\\\"\\\"}g7a6a@a\\\"\\\",2):f(\\\"\\\"{g:a?aMbKaKa6a?e:a@aEa2a|gZfMbbgki>a:b1a-gemUf\\\"\\\",2):f(\\\"\\\"{bHa4atcDiGB0j>Y0jBU\\\"\\\",2):f(\\\"\\\"}bJaMa\\\"\\\",2):f(\\\"\\\"}bUb0j|?JaJaUa-bJaMdJa8bY*;a8bNrKa8bNr/S0j\\\"\\\",2):f(\\\"\\\"}bT17tGB9bKaK62,TaK"));
$write("%s",("6K6tQGB3:JaLaJa8bXJGBd4coa8bNa4uGB:b+b>Y~4aka\\\"\\\",2):f(\\\"\\\"}bJaHaJa8b93a/aHaJaJaJYVa;aK6Ua:aUa:aY*uiSfQfFl4aX/sbsb2be3^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'mauiDa-a;C*b-a<6asa;,Ue>a4j\\\"\\\",2):f(\\\"\\\"{gKaKa|gZfx6cgaagPjkg|6esasbvh*b-a/bxcHa|fCke3c8c\\\"\\\",2):f(\\\"\\\"}b\\\"\\\",2):f(\\\"\\\"{gph\\\"\\\",2):f(\\\"\\\"{gvg1a-g\\\"\\\",2):f(\\\"\\\"{bHaCkRf-e:a:a\\\"\\\",2):f(\\\"\\\"}bHa?a\\\"\\\",2):f(\\\"\\\"{gJa\\\"\\\",2):f(\\\"\\\"}b5aAdte@a1a-g/iCkxcpb7anb2b:b\\\"\\\",2):f(\\\"\\\"{g2f?j@d-aIfdkxcHa>a1a-gigggsi-aUf/iwiRf-f-gSf|fCkzeSgwiHabk;a/aCh<b+hVh<apb/aChVhnb<a<a7b:b\\\"\\\",2):f(\\\"\\\"{g/aCh-f-g+gFa+i|b1aki3b:b\\\"\\\",2):f(\\\"\\\"{gJa7bH"));
$write("%s",("aCkHaUe,iCe|bxc3b0a:b\\\"\\\",2):f(\\\"\\\"{gIa|bzeJa|k5buaQbwi<b=a-a<m*c3bxdUem3aea|b9ai3edb2bMa7apb4Vphnhlhjh9apbqhohmhkhKcdc/bPcgfvfNhIh7a4V/k-kMa<m*cEc,dJa>a2aIfyjMgMa<m|b;i+cai6a/3iUaxd/Z8g/aCh=aoiRaTtCdTtkbG,ZUoiZj6a7b5abkRfwb|jUe2b5a9gXiD@hcZrNiNiPu0c/bxd;a;hnj%?aea6a2bJ>esc*B4R6a\\\"\\\",2):f(\\\"\\\"}n2a5a.l@J\\\"\\\",2):f(\\\"\\\"}g6hik>@Ni6aThjnHa1dmdKhRfVkKkHa:eVkKk/l<b3bxd6aHh7kOhmd+Kjijixb8iacPa;a,bNh2xfbpbubld1bZb-Fnbpgtjrjhi5YQiUkuhSk3j<b<b<bEj:b;j<b<b,cJjGjNqJjEa:k\\\"\\\",2):f(\\\"\\\"}k,cBjLi9a7b6g-aht,b,cJj=a9aULxbq3e13ecaBj13iC3a13ifaJb7bdS3fkacdaG>a9a</)3blaFqkoj6k,cJji3asadmhh.bfh,cJjsbHa\\\"\\\",2):f(\\\"\\\"}gu5ciaUjCjCaKi:6aka6jgk3j<bze;Cc/3gda1k3m3fvb;kKi6a<bjibjgp*Z0Rd12a2aAHdkNk/iwb|jRf@a>anc:e7b5aWf=aKcU4uk5a,bJa6a-bJaJaubJa7b5aUgwb|jHa:e-b9a9b9a1kdkyg>am3aya01dkyg"));
$write("%s",("@a>a:a|b9a0b9a@a>aBBa?a>e|bPg9bJa0bdkyg-b9a1k9aCaAaJa9bdknbJa6a|b5a,bRf:e-b/kW3-aO;a(azi*Z0RuiAHyg8bAdFh-aAH*b.bbb-aAHyg7u3jlbAHKc=ie\\\"\\\",2):f(\\\"\\\"{xd6a-b9a8b9a7bJcJayb>aduji>aJa*c@dxc?b,bg:>aJa-b=lteUe@a>a<a2b5aDcP9:atcJaubKdZ\\\"\\\",2):f(\\\"\\\"}5Y,bD@JaUgq7eeaIkGks;e)cRkPkpb;awb|jrls\\\"\\\",2):f(\\\"\\\"{.B\\\"\\\",2):f(\\\"\\\"}Z4T4PBJ6F\\\"\\\",2):f(\\\"\\\"{ZJdHdtlzn=n7lam-n+n@nBn@a=nJlF|3|mbM5\\\"\\\",2):f(\\\"\\\"{bC0<V1b-xTab67rb6\\\"\\\",2):f(\\\"\\\"{Y?EW6/bZTt*xWEalsp,-X0bV<aGEaUvv.r9Ea37y=GWuV:q/b03co:p\\\"\\\",2):f(\\\"\\\"}N\\\"\\\",2):f(\\\"\\\"}K,olh=aq9L|PaDJub6wFOM,q>Ta2br38bYahbjbvbDu?aupibDajb<pU-/8lb6bu8y@k5a$d9AE7<RBaa.|bW6=/g=ebGxt04@:zDpRoB=A0Fr3Smbp,TafbIo3\\\"\\\",2):f(\\\"\\\"{X|:y/IqyYambn<;qTooNt.XL5bMwvozLOqv8Zx4shbRaDa1Q\\\"\\\",2):f(\\\"\\\"{6YaglK?p:4|b-/5lboYc.RDEKl.q\\\"\\\",2):f(\\\"\\\"}6rPaYAyDuu\\\"\\\""));
$write("%s",(",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"}eFBaJQ@t?BvbKyib+b-2YtcxF|dbPa@RjbvbLtnB\\\"\\\",2):f(\\\"\\\"{bWaFas6GxjbXhkbiP6\\\"\\\",2):f(\\\"\\\"}@EAs1E<a03Ypo4ruXa9B>qUP\\\"\\\",2):f(\\\"\\\"}FaQA*@XY+kb2o+x2bRa*xw=k|tU>as:U@VaufYhZaDj6uHuy:?eubEu3yQa-Vv=5s*6czd5oFzz8spZavONVUyZ+Z:XFpS-1ZpG*HwSaau+;cbDa*b<aJAfg0IXGN6\\\"\\\",2):f(\\\"\\\"{bWaO1gbXaQtBaLTVaZ|k|uu.K2qGR2|4|BKaz.bVtZuPER*Ckwwg.YR,p3s@aR|QoUC6b+bYaFa/AA@kb@ta\\\"\\\",2):f(\\\"\\\"{fb7q-bInPa,bxh2qInnFEnVnO,i>6wFO+bG/;*?a9|+bG/Nj03vx>aYaWE97lbzsT3>:*srxc|gCjiuXrxkoio-8pog\\\"\\\",2):f(\\\"\\\"{oUlo*7uAXPK+=OInx-mbpo|XOrApjbQFK/N|dx;oRTPTNTkhWaJT$6c\\\"\\\",2):f(\\\"\\\"}a0<poJxET?aPXQXC/?Tdo*bpoEGE,Y3akcdb7ojbVa@aib0<jbzsfb?:Lz-6D;5tPp0<c;fob6lbpoyx1Q4bkh,NUZgbyx1QCiN8mbAv+4RaTAOSL-Pr,bb6zr4V;v|5Ra,b09.,N|0<1VAvEav4y\\\"\\\",2):f(\\\"\\\"{@Sb6L0i|e0*vWnvb=ymb9bdbWn6bAvEa"));
$write("%s",("vbXIPpNBc;<p+SWn25BaEacbAvEaFRWn-6UaQ3aEa+RstcovOZp>a-0O6c;GKPaV|09K/-btqjb7\\\"\\\",2):f(\\\"\\\"{A2gbyx\\\"\\\",2):f(\\\"\\\"}5kbA2WQrsdoHyDajbksN;&6cJbHyDaOq4pTB1b3<ULSxdo..-Q3x7bNQHhX-1jDaQ-FO00;6L1\\\"\\\",2):f(\\\"\\\"{bc3=a1bu\\\"\\\",2):f(\\\"\\\"}?eRMDxDa-o,bXP3hpRabnRmblR9\\\"\\\",2):f(\\\"\\\"}DafhFOn.M*hb?Cq1p>dbq>;6Qa?a,b1Q:k,blb3b+psp;6WQqLv0GpxM<tq>;6b+jbebXs\\\"\\\",2):f(\\\"\\\"}3e.blb=TtpyhCpWagx6p,\\\"\\\",2):f(\\\"\\\"}hbRaqxq>;6Mn<aDaWQ/u?;Ta/Fhwnm0bubBakb|o\\\"\\\",2):f(\\\"\\\"{zhmV3gbGotbINhbfbtb=a2E7=pOT>Zpj-F;zbLvsqRot0XBlb>a?p/8K0cIlb-JPT<Blb,6c~b<3<3<30Vmb\\\"\\\",2):f(\\\"\\\"{bQtZ=0|vb=a44FsNlc\\\"\\\",2):f(\\\"\\\"{hbb+iblhc3Z06\\\"\\\",2):f(\\\"\\\"}44mb\\\"\\\",2):f(\\\"\\\"{bE0C@W=hb@B*b;kCp6Z*bDa;6YY=aDaW20-6btb\\\"\\\",2):f(\\\"\\\"}-2:44lslhCwdz*<TaZ:IrzyEan\\\"\\\",2):f(\\\"\\\"}|4aRb>Ez67|O2gbOaLps4n8gbdL7|7bm\\\"\\\",2):f(\\\"\\\"}C?"));
$write("%s",("RCV-4bE46Am81;iQBXUpg2g8m81;:=q0l7v,Bt9P5@ub*=OaCG61K0jbujTafb?a:y\\\"\\\",2):f(\\\"\\\"{*mb2|+bE0:4+yVFe,t0Pa>ykbLqB?4G,pFu/b6o3ZvrmvVFZ:blPS4bN*AqXK<qwb?a:@eydyp|sPtWOPS4yPolN8-2=k9-+iXzs6beo5EYV0bBE7CwQ9fPaUaoEXaaw39QB;,YV/,e32bH624Q-3hLp2bWa.b|wwzQvxbWayb0bdN2b;+lU<WTEusTanCwjQaoP0-?p>a4bhJ.kr2nFTtDzXaW71*-hMWBaGapMMvpE2bTA:36/9wo8tUFa|pyFH\\\"\\\",2):f(\\\"\\\"}eN2oNl2u0bCajbH+/bdx6bz.Ta6*iscW=EsRe\\\"\\\",2):f(\\\"\\\"{BKa=mvCavlTa3b8DI*A3JAXaX+/|dSsu:sybw;o8tU4b7b9rK\\\"\\\",2):f(\\\"\\\"{yb,2xb,Xvu>&6d&dAvRslW3,k+<r:r8r6rd+55ZEN*5|\\\"\\\",2):f(\\\"\\\"}bKCM>xrRa6*2bTA=|cbNVTooV3b?Peb\\\"\\\",2):f(\\\"\\\"{2Cakb\\\"\\\",2):f(\\\"\\\"{v*R@EOt?pmb+\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"{bbb\\\"\\\",2):f(\\\"\\\"{qjYzb:3y\\\"\\\",2):f(\\\"\\\"}p;v\\\"\\\",2):f(\\\"\\\"}t\\\"\\\",2):f(\\\"\\\"}r\\\"\\\",2):f(\\\"\\\"}Hr:yTEjLnx@.XH5o=Xe6K/uF1*5obViN/G0bXa"));
$write("%s",("hb\\\"\\\",2):f(\\\"\\\"{bG/Waqw7-E\\\"\\\",2):f(\\\"\\\"}XHkqfbnK*b,n4b5b9bcqYaSxUa:7B?\\\"\\\",2):f(\\\"\\\"{rntZq+b|p?a9b0bRpzbqsyb1v3baBGV5byp.kc<ScSa+v:*ZLib0bv5?253Ra?;9<Ba5of3lWXa1;+bhmjiAT7,GB;YBE9*CavJhb-bC,U6:9,6cIao0E*VaX96,|beb>yX9fhF*:tTaF7N**;xxLs<aUaHSXh5o8-Xw=|>aGB8.T0VCmVibd*^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'3a*cRaNaJx@Y7,*bS*SG;,?YNa*by,2J3<cb-r-6oDY\\\"\\\",2):f(\\\"\\\"{c6r6Z02|K*qxC=9bkbn*Gaf:K1ib7*PrUaToVC;sIIy.Uy\\\"\\\",2):f(\\\"\\\"}br2h6/,cz,b97\\\"\\\",2):f(\\\"\\\"{*t-\\\"\\\",2):f(\\\"\\\"{7hq=|nvlvjv>@G@XBg00\\\"\\\",2):f(\\\"\\\"{3b*9yb+rgw4xq2KVaq1x,tawQ4/bmtZaryzzJ>avOnEae3Awg0a,6\\\"\\\",2):f(\\\"\\\"}M.+b"));
$write("%s",("yQ|b6\\\"\\\",2):f(\\\"\\\"}01vBM.fb1AZaJ\\\"\\\",2):f(\\\"\\\"{@aiOoEPM9d\\\"\\\",2):f(\\\"\\\"}dTo1bUy*w9b6L5@8b8p\\\"\\\",2):f(\\\"\\\"}G8>C.1bBXf?9=|b|vXQBaiz8BXs\\\"\\\",2):f(\\\"\\\"{sd,?u5vEaV4cb\\\\\\\"\\\"),\\\\n(\\\\\\\"\\\"Aa26ubDZubb,cGabi|6bm+?a6vV4cbKIUy25ibfwU6\\\"\\\",2):f(\\\"\\\"{2=YPaFRhT=ZcGab.bczzbVao;PzubEantJz*zRM7bVB:+5<+Rm>?hnwDiyz9,R6KUC|r2p2db5<rPau@zL\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"{tN0H,TD-Q-0|bTamvkv3b,\\\"\\\",2):f(\\\"\\\"}ZMrS+79zO9\\\"\\\",2):f(\\\"\\\"{r8zTUfq=z6b<acbX?vpPa26Xilb;,YVPahTypupFRkbh2jbb0TBCGDJ=quFyvFIlW-b\\\"\\\",2):f(\\\"\\\"}zNdea@,O9l4aXbF+q+z;.bCSt4K3p3;-Wa9Ta@9q0v7b3bU+,53baIJ9Za9bfb9SE0fbs;jb?v0blG\\\"\\\",2):f(\\\"\\\"{*t-Ua|PC0W;QakK<E/bxhy?ibww5J1b>R\\\"\\\",2):f(\\\"\\\"{bG/+j:UQarr:7Wa5oGBAxnk0rdIYt7bVp,b3x<I58=|Ea6GUa-qXpLn6BQaDrNlfbRaUz?az8atbmt3r:5M.h>/-?vd<l,j,4bi6K\\\"\\\",2):f(\\\"\\\"{wb?aYs3bn8CC?=U"));
$write("%s",("Zt6;v+x\\\"\\\",2):f(\\\"\\\"}by;QVg29P8-Oa=Eor4Msuwb7umtcbDa7\\\"\\\",2):f(\\\"\\\"{?a1hlT@EubabDwNaX|N8kbC7*6c)d|uubebcbDa0u4|KyJTab\\\"\\\",2):f(\\\"\\\"{0fyU8Paotupu6s6qyvb*b1=@z>zQ4AaTDhyvGybv7vb4Cd*Mv.TKINr/bB1zyks=ZXaZ2;<ty7U9R?a\\\"\\\",2):f(\\\"\\\"{O/b7>+JA,vbc4\\\"\\\",2):f(\\\"\\\"{2*rmGZ-A,ibn:LK.q6,+5yb/zFa-Ukb:yKhE*Y9Fa8bqo@|JyCaUa3/*b=Me<\\\"\\\",2):f(\\\"\\\"{8Lu7bb<.b2.><4yZaQaJ-bbr@h,\\\"\\\",2):f(\\\"\\\"}s/-\\\"\\\",2):f(\\\"\\\"{bbb2E\\\"\\\",2):f(\\\"\\\"}GWaZano-umbBf1VWaBaNht,gbXan7+vAae0i|.b<m@zGapMJ=bAmb*q;vQa|Ehw5v+uerfWo9xbNacJ,vW%=dfbf?+vAa7vybr6A7AaJvXBWynLc66bqT9zub+:Na<IabTieSfbcIlb5vgbp:XaAau7hom\\\"\\\",2):f(\\\"\\\"}Yac;e=VV4VpGvX?iG/RXmbUA>Da|cp5Cawj9bjb1bNyCa\\\"\\\",2):f(\\\"\\\"{buMMBGUGaf:RwaDG4\\\"\\\",2):f(\\\"\\\"{bc4kb>tSpLvMB/xkb<V+5<IDr++G/LvQ*eFXaGa?YjAgbQ3ubnsFazb@>8b8bQaFaXin1S,>tw=GapMvb>aL.vb>aPaTo"));
$write("%s",("212bVC||\\\"\\\",2):f(\\\"\\\"{0PaFnupIzPn|Ifm9<BauqU1MXM*X4?aYUPz6v<uNj0b..;qWaRaDOa.|bdL*C25f4NdCaibBCUa2g0-uk2hkbJFJ.9-3b/br,v/5|LK?\\\"\\\",2):f(\\\"\\\"{UaOqJ3>a=itrdYQaK33x|bTaw;^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'3cu3a-cPat->PC1+@4b5|cPK3Pa,p<w\\\"\\\",2):f(\\\"\\\"}EUw7,7CUa>aK3PaC1ubcb\\\"\\\",2):f(\\\"\\\"{v>aPa78D/lX+x++FqFg2bVBqv+<\\\"\\\",2):f(\\\"\\\"}bhb?a4WWaNr5wvAcbjx.\\\"\\\",2):f(\\\"\\\"}lLDX5oVXKy8sn\\\"\\\",2):f(\\\"\\\"}f.Vp3svJU6?a?:M.e=L1wsQ*BOCayb-Hh+Is4bX5i9f\\\"\\\",2):f(\\\"\\\"}sM8JmoX+UaEq<aS3/8abNEh,\\\"\\\",2):f(\\\"\\\"{fT*hJWBDa;<Raxbyb0rKS.b6??vUytRevhs*6ekacb?Bg:>U=a/3a>bVuQo+vybR8/-avvqYAMqs;+oxb.b\\\"\\\",2"));
$write("%s",("):f(\\\"\\\"}F31gw5b8qjiGW>vAy-oKrVnC2iA<a\\\"\\\",2):f(\\\"\\\"{7Wa<L/PA00hVv8q1V+*29?5RDX\\\"\\\",2):f(\\\"\\\"{yU0hVP>aubFaB|evosN95o6v2q57tqqr+J1bO\\\"\\\",2):f(\\\"\\\"{KUKSlbn:@0UajiPScZ40q3e~b:/+7TDxW,qE|Fa5byx+rE+db|bxyDM+:5b0rJYfB/b:3xx*vlwpW,blbs9E|XlC7zNtb:3g>o4l7CRQT-+Dyh\\\"\\\",2):f(\\\"\\\"{6fqTXacJA*Hv+bIvFDUAwbnhd\\\"\\\",2):f(\\\"\\\"{2rfx$6cbbexdK<Yfx/bNUEafbf?.bPa.d,vWPWy<,<aOW\\\"\\\",2):f(\\\"\\\"}zsM\\\"\\\",2):f(\\\"\\\"}zuuH0vb4CFa/b/bcGU3?u.I?;d|tO/bY6F@+bPnNaOUdK\\\"\\\",2):f(\\\"\\\"{yU3aca4qS3amcVz6@ey|pVp-b5rT**\\\"\\\",2):f(\\\"\\\"}fvJ4d,mvkvUCJZ5bp1X>E+-6UamG7yPXakYsybBa5om5:4i-\\\"\\\",2):f(\\\"\\\"}ztbU,srzbJv+be+BaZaoCJ?zv<L.b0IoA6|8DBXkA1JQFBauv=T:UttE*l+1V4;2siAFacJvvvf1b;\\\"\\\",2):f(\\\"\\\"}7yjiPSp:X\\\"\\\",2):f(\\\"\\\"}<aQ/2b7blS/bxhjiuXT3@XwbvvzVO+&6cvd7gujlb.H2vS,,b?h;*DFebp:<E,Y\\\"\\\",2):f(\\\"\\\"{b>ryFOXxvOavv"));
$write("%s",("tvNl2u|paD.4D8-bYR?5RDW7TIPqiba@i-M7dGGakwM?/b9<7vld?uNa@udNjry,Mzyb93H?P9Fs93jbKSBa=tP9Fsz;+\\\"\\\",2):f(\\\"\\\"{qUfb?aIGdz=u8bVa2;<aK\\\"\\\",2):f(\\\"\\\"{wN8BPyybAawjzM?a8b/b5tPI5bCaoEr2M\\\"\\\",2):f(\\\"\\\"{Vaw+is4@fh5bhhablNFO0jN=6;4;OaZa3gPI5b7bp:GYp,Mo.;Van80|8-c2q07<2x?aKo8HpR4b0-Y<YVa;hr4bFq|6csd0bg=EGnC,AixZs/bn=++Fq1:FqFzcxLunvQvAw?Fp,BKa=abFMW<f5\\\"\\\",2):f(\\\"\\\"{u,blblvF:B@WaJTy.m60-Uo;q@aYg<ExW,yTp:Qn75<HKn<3b;:QaSay.c?ji7,0s7ST<Zx+x7CK?O,*=*wjr*4xJ1*lSs4Fqzbzb4bQaFo|IOajb+x7bS|+d+j1JoG>Z8M2bZanCdbk0/bk+?C4p4b+x7C<|B=O.GKkb<s9bn=c?UYA*tQQK9b.@x3HNT0DaNamoBWQ33U3,kb*bUFoosrkbZ61;/qrz6d\\\"\\\",2):f(\\\"\\\"{Ek2a751b9B?@v.\\\"\\\",2):f(\\\"\\\"}bgb|X.xI+x.jok..s<aSad<.KFa>?^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^32^[2fha\\\"\\\",2):f(\\\"\\"));
$write("%s",("\"})1(f\\\"\\\",2):f(\\\"\\\"{#v3mja51(f\\\"\\\",2):f(\\\"\\\"{#,4353(za199(f\\\"\\\",2):f(\\\"\\\"{#(ntnirpn\\\"\\\",2):f(\\\"\\\"})215(f\\\"\\\",2):f(\\\"\\\"{#)|4[|4aUc.s:YQaSa7-x8o@Fa>?5oj@Di4bzbRD4bVa?E/tyv>aTVm@/t.bD,>qVaGaYMvbEajO094GB.d</bcGL|swbb>awbDplbx3Sak.3wu@fAybq0g4l.4bAaibDa|8a2BqJ-3b0<FIkso.dbHn?aD,Rr*bt@*boU,dEaH,>qVautk|lbf54bEa3b\\\"\\\",2):f(\\\"\\\"}5ZQ@ab.T8J+KIc<y\\\"\\\",2):f(\\\"\\\"{tbEr5t7Ct-VaaU=<S|/bAte3cDak\\\"\\\",2):f(\\\"\\\"}b+bs/XaMvK0/rhbD-Yau|jb2EtQi9c+dh+uof3UaoE,ySyt9Za;6oNEYCa?agx+K\\\"\\\",2):f(\\\"\\\"}b5o8p-UWaubTa>ZQvJo7\\\"\\\",2):f(\\\"\\\"{q,-C@rUBNargeLD,BV*4<aSaUA@rI*+bZaYJ*9UyAB5<y.-bctZbkrnu\\\"\\\",2):f(\\\"\\\"}qDaU-ABebGaYVUV+yzbT,xb=aVa@;S,hTjdtrjbwbF;O;q:|pa;EauVR6c24M*bCC\\\"\\\",2):f(\\\"\\\"{bzp<aRaebhbmbRv\\\"\\\",2):f(\\\"\\\"}beo>VEa-FqWQ3mqsV+bX:-t0b3UT,6bQavb0p3|1vMXZsN|jb9b2bRaWa=<Hw.bl2t,zG+b"));
$write("%s",("HH5Ih+><fvq7OrQD.b::c<..wwTa9b1seb*fJdRb|vm\\\"\\\",2):f(\\\"\\\"}0*TaX\\\"\\\",2):f(\\\"\\\"{/A1pMvP6Baw=eB02xW8DhLkbDa><qQh+Qab.BVS|Na9BS*T>y1abf?Ua5wg,r,BV7bybNa*b9bWotqn:.bbYX-Va9ow.gbv5M\\\"\\\",2):f(\\\"\\\"{a5t9srK43wR:ybMpwUJy:/Ya.x8zMq8D1bN;3b4-m6;*t+e0uzpSXOr-hHa:b<3QaC0K*IhhLkb3UCG5:C,6bb<1x;++rgwf4?ag4U4|bj5JQ5s3se3.Ezb,ETyuEqoD+wbD//LoEgb2E4s,b\\\"\\\",2):f(\\\"\\\"}0spYy9X=tVoOp,VX\\\"\\\",2):f(\\\"\\\"{oAbbebJYab2Es\\\"\\\",2):f(\\\"\\\"{.B\\\"\\\",2):f(\\\"\\\"}Z.l@Jy@BJ3RR.\\\"\\\",2):f(\\\"\\\"{bS,YnW39UghdwuAUmbl0L|/G-4qqlb|rwZE4CIZW>r|w-sCs1vBuToQaldUadb9<<E*bOXHSXaXV3sJv.bKUj5xh5Z,vNzr\\\"\\\",2):f(\\\"\\\"}p>QSeTwbjJ-bLs@aYaJYwX\\\"\\\",2):f(\\\"\\\"}bm\\\"\\\",2):f(\\\"\\\"}g2Z*fbg7O647yxd7mbKqWQTa-bwb0bmbqwp:q;o;,p3bW\\\"\\\",2):f(\\\"\\\"}U=JF?;Kv<a9<+:\\\"\\\",2):f(\\\"\\\"}swbdbPthH,S<aPa\\\"\\\",2):f(\\\"\\\"{lCud|0b\\\"\\\",2):f(\\\"\\\"}E,pmh<"));
$write("%s",("a5oX<TsBuRv;*3b0bXaa;,SM|-b-6/P<a,bn>U,hb,\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}bsqF@ntBaOS<CvpA=RvBZ0p&6a#c0D*Z0RMuldureocbfbjbttK0nK*bIHkrtJZq+b|p?a9b0bRpG458962bibfP7oVyCqOHMH4xMp.IVJd|.byzibGXC@\\\"\\\",2):f(\\\"\\\"}-2<WaLqZa7td|.bPakS@auq<aQ/::T8-6bbm1Voe,uxp3kbPq?25om60b;\\\"\\\",2):f(\\\"\\\"{?aNj9E<|=a/b..@0pql;PnTa4vQDQqr>ebK0T9Zs9pcJuxQaZ+SGdvA3gTaMTj9*uxb.b\\\"\\\",2):f(\\\"\\\"}boUA77*TBjbF27b<MlbTaJ6,o/G/bwyMIG;t6uJ96SGhoxbybHH8H/,ibE\\\"\\\",2):f(\\\"\\\"{cx7CWaN|2\\\"\\\",2):f(\\\"\\\"}=d(df\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{:\\\"\\\",2):f(\\\"\\\"}@8D\\\"\\\",2):f(\\\"\\\"{M9b5b\\\"\\\",2):f(\\\"\\\"}b+bAoub.b4*Xi.Z@ryLWzp,8b2wE*@acGM|n:JSQa4Gzslb4b;rVJO:LuXo47f-GBVabbRa*>LrW2DaN;+bLrCk7v<awb7vMIBaD+zFb3|8gvqrDOd@CwJ.|blbubD-J\\\"\\\",2):f(\\\"\\\"}fb4|0hC-Ba>=N.46VaAqwbnsKDJ.jOYJKDVaqBEazVHR@acbj57v9bksfbg<r\\\"\\\",2):f(\\\"\\"));
$write("%s",("\"}*>Lrfo4|xbfvfb:JE0:J0bBZD-N;+b4|*>Lr.dYh9<r\\\"\\\",2):f(\\\"\\\"}*>GucJqr@a\\\"\\\",2):f(\\\"\\\"{uQa@a+bh6UF<|KDlbHK0bjbHK0bn7=a/5B=.6coajbC;5bf-K\\\"\\\",2):f(\\\"\\\"{w4|fc3imaxbZ2*dybPa9ge3aIckbjbubO:C\\\"\\\",2):f(\\\"\\\"}.Q6Uckjx9b*\\\"\\\",2):f(\\\"\\\"{qB**-b.Kp3?5M.Xo8t5gE6yOn=4:Yaw9<Er>tbokbb?akY\\\"\\\",2):f(\\\"\\\"{b@|9b1sZq\\\"\\\",2):f(\\\"\\\"{*|898wUmA;KX=.+i,.wJv@a?hcbRPjidBXa9fPaeQbbtqi,Yne0ctrgX@xFm|A=xbU=VvAa/55tcxC;<E@MU/+b|X=u2bn08bNJE*4u2x*;|8Gxjbm|fm+bv/Pay*dJ=ahTLvTa2ht@Lp\\\"\\\",2):f(\\\"\\\"{bG/9B<Y5bAaLvS14pcvQE&6cpdp@2.5bH+aT\\\"\\\",2):f(\\\"\\\"}zdVZ0Zy/-:,MqHtjiPSkb1pjb5bAan,8D|:J309aw-bdV*=fbnKL|jiH\\\"\\\",2):f(\\\"\\\"{b?o*drx6;?|:E0TD=aX|R5Iy?FU+I+H0?ac131VU<awbA*:D+\\\"\\\",2):f(\\\"\\\"}z;f+FNw=4Bso\\\"\\\",2):f(\\\"\\\"{LdFDa4sBSMtW,6bn>3smGkZ\\\"\\\",2):f(\\\"\\\"{?RaR5sM=Q-VfvHS,b4AB.yIGwMvULH?:Dabi0vqB.yIZs6bV"));
$write("%s",("<E7s1f8abWPmb2|ibTtjbb0,b<an:fbEa7-pGvXzygMiXzb9v6rJ\\\"\\\",2):f(\\\"\\\"{C=VoJA.blSUQjbsoXaatv6cOcYs6teu-QZ+3baO@RybRaDJybHKU?Za6-7\\\"\\\",2):f(\\\"\\\"{Tomq3wmJR*Fs5Jmo9v6r1:<YnoJr2bMo/byb5oXafx98/A9bJ0hb@zujB|Bu5o/I.bv7iO9b:10zb*l7@?zb>aczJpn,f5s*6b1,r=6b;6TZkb:t/-8b:Y=?9g*b;F9AyVZagQDpjbp3kbmtyOQa/bTaAo=K\\\"\\\",2):f(\\\"\\\"}JQ-FOOTF|ZaX\\\"\\\",2):f(\\\"\\\"{gov7,iH6gbLs:zLs0tE2mbZa0j0bmbUygxKrl>kFL1Vt)Ua-auoxbdb+b\\\"\\\",2):f(\\\"\\\"{bur37W-ab,bcx:+UM,q9b5;Xy50<YI:,6cCaubebt+au06?aPX4MoDabay1-au8p5<4ufbtb.bT*P|>SiuM4Dj>aZUETubZagR?3a)aabO-PXp:oDdMFp;DWTO:aNgbm\\\"\\\",2):f(\\\"\\\"}g215k5ETO1/3akaeH/1-1uy+4g3aY2\\\"\\\",2):f(\\\"\\\"{bk\\\"\\\",2):f(\\\"\\\"}+b0-uyydZanC=HZOu|JhVayb1v2hX\\\"\\\",2):f(\\\"\\\"{jqG*iuL=tQZ@oE/b3xZxPzBSmGntyK-bE0bb+pG2e0zv/7fvUA/b\\\"\\\",2):f(\\\"\\\"}zNz.x/4k@PqJqfbzbE6/z8Zwb@ah+Bsaoac/5Fz"));
$write("%s",("D,2=@Yn+orqLpj6Ygw>B094lt<1X,B/XTpGaxTfv8|-1Pqor/zW*OWvO3|LnYYe0.Aabq08=:p8-QxoNWa8;,7lbCaPP/52qKY3bkP/9CaXl<ox3oCQ/+b<aFar6sM\\\"\\\",2):f(\\\"\\\"{b=aubUVxWjiV;+b>afbF|Va|v5n@,vb?a*95oW3k>xI5bGvgc=v.7mAB7D3Q*Vz\\\"\\\",2):f(\\\"\\\"}JL1W5HvY*<|e0e\\\"\\\",2):f(\\\"\\\"}W5**UafxzF;vfbkbdI3b1Jv8ouo\\\"\\\",2):f(\\\"\\\"},*jb9JUpvUmWq0P6-0U=\\\"\\\",2):f(\\\"\\\"}J=|GaCTkb@P\\\"\\\",2):f(\\\"\\\"{bHN5bwsirpGbbzpUx\\\"\\\",2):f(\\\"\\\"}bk0dbi\\\"\\\",2):f(\\\"\\\"}6b5bxGzbQkCiG4ybNsB3Y*\\\"\\\",2):f(\\\"\\\"}8/51l5R3PE56V,bibsMHvzQIG3b7/l,xbt\\\"\\\",2):f(\\\"\\\"}4b5owb\\\"\\\",2):f(\\\"\\\"}C@O*rk,wbyLItcGzb2bbr\\\"\\\",2):f(\\\"\\\"}bL|irSa+\\\"\\\",2):f(\\\"\\\"{.5I:Ksfqyb29Ca0TP-+PJVvv/8d..b.bQ9lb41Swgrr6eB|bEa5b1JI,kqf5w.nt>p<a75ox-4ws\\\"\\\",2):f(\\\"\\\"}VlbB62qDngb;C1bC\\\"\\\",2):f(\\\"\\\"{Jh0qgwR?MqLKQ9mCEUS*9=Ba4Gzbk+uy1;m|k|ZafqFp/SgbeDk|iynu/GoNJh|s8T1TebF1,"));
$write("%s",("\\\"\\\",2):f(\\\"\\\"{bbn:m\\\"\\\",2):f(\\\"\\\"}wbfbXsNN0VH?+r,b@8.dPa/Eg=vx0bji=5StN=Dap6JxLpR?21/bdwy@B55Ty@3TEa|b|PGaEShbCuJ=kbZa6t?aBaJFeVSa9bWTk|xl1bQH5/xbLDPaUAR|1*dc9TfcSa1ss9,pmS6b:UMEG@Na6b7qe=Q*nsab@a.5U8:phyv94t2|kbgvI+;Kz.i>lbG/1A3bOa.kG/ubZhVvl4tbp3;,0,bbG\\\"\\\",2):f(\\\"\\\"}/,5ox6Y\\\"\\\",2):f(\\\"\\\"{E|jbm\\\"\\\",2):f(\\\"\\\"}Ragrqu<te=97InS*\\\"\\\",2):f(\\\"\\\"{bhU5bQaU4zb|O\\\"\\\",2):f(\\\"\\\"{bPafBRaPaI:>pE|*5lb97Sai97CTaE,MyVakbuNffRtgr,\\\"\\\",2):f(\\\"\\\"}Njk0Qtkbwb1bZ:EyWa=aSaVaR8x\\\"\\\",2):f(\\\"\\\"{C,hb1,2y<|jirCbozyXaD4utE,8b|bU.\\\"\\\",2):f(\\\"\\\"{3-BU.1Ptb/p3bMBTab.2batlbixr?/12\\\"\\\",2):f(\\\"\\\"}m*0\\\"\\\",2):f(\\\"\\\"}-0o@j5Dn>twS0b>akb2h5gkb3wk2URYaLs0I-bDaR|Sa0b95Sahw/vVCHSPEuz.K5oebEa1wXJW6,bzbaoTayPjiCrwSv4SaN|xx3SubWog*F0wsQa2E8b-bORj:5b-bvOXJTa53*wEad31bQE9P;KJy7>Nap6FRMLsseBkb|PQatjp65b"));
$write("%s",("vbYaRrhbo;Jy7/\\\"\\\",2):f(\\\"\\\"}bUapEks53aoybtb\\\"\\\",2):f(\\\"\\\"{P>RY|6+Na-2.uerIn?u\\\"\\\",2):f(\\\"\\\"{bDnLtXFyJAa\\\"\\\",2):f(\\\"\\\"{bdbFaZ/CaQBFIhb\\\"\\\",2):f(\\\"\\\"}zfbjd=aIz6?/9ab2hy@1R7F2Pw>G57N5NH6uHP22bCacbyLbb-8M\\\"\\\",2):f(\\\"\\\"{+1-/:qfv*b+bPavy*bv7BxIrW|bRfhYaQH>qe/@9W|QacxVa9byAgbjbyADa@Fo72b9o*?>q0pyAe\\\"\\\",2):f(\\\"\\\"}Qt,b4y>@WmtzX@7sc41Qk|fyhxkA.3/AhxPak5jis5K6Oa*o2brqDa<qOauy?aQok6bAiJ<trPQaWao\\\"\\\",2):f(\\\"\\\"}BtnChw8bh+UaAa:4TtIo/Noobb4B6bkbhb?v|\\\"\\\",2):f(\\\"\\\"{QaSOm\\\"\\\",2):f(\\\"\\\"}ub+/<thbE6cbTanKaqEa\\\"\\\",2):f(\\\"\\\"{qp>\\\"\\\",2):f(\\\"\\\"{q3v7vbE|bA=@>ls6fhlDxR|KGEqL3kbDqcbN|DnDad7abi\\\"\\\",2):f(\\\"\\\"}Datqs\\\"\\\",2):f(\\\"\\\"{8NT.r<6N=wubRrO1ErILIsAtabBaU/cbZ7xb?y9p,A8b2bS3nF15W-|zdx8b\\\"\\\",2):f(\\\"\\\"}5OaA16bGuaA5<QaauY\\\"\\\",2):f(\\\"\\\"{EaD\\\"\\\",2):f(\\\"\\\"{4bjih*.\\\"\\\",2):f(\\\"\\\"}2bbbi\\\"\\\""));
$write("%s",(",2):f(\\\"\\\"}7\\\"\\\",2):f(\\\"\\\"}ub1b-hB6nsw9*w2K<zYadb1w/buz0bvF6bhxPslb6uHJF*aD7q3/TD4H-:/bQaUajbMB0g8bRrYqybxMSaQa753bN|fqfbX@<abbQnZKfb25-4PDnhj9FaYaQ3+bwxEaVyn:-1Sae0Z=yq+7F**4\\\"\\\",2):f(\\\"\\\"{qVC@*/EwjO4db3:ibS-5b0b2b7>WaV=Zh*bF=b<T9@u.NdbXBMGX@Pu8F1D?L4bLsbbMqcrg2/bt9\\\"\\\",2):f(\\\"\\\"{?9b1-+:7bMh;Khb5E+FZ01t?a4C>a\\\"\\\",2):f(\\\"\\\"{9R*foXaIse3Wa\\\"\\\",2):f(\\\"\\\"{wD4lbJ9brBKydjbX@;?5qjiEM2?S5YaV3>qXB\\\"\\\",2):f(\\\"\\\"}burW,,=B\\\"\\\",2):f(\\\"\\\"}abxM9bu\\\"\\\",2):f(\\\"\\\"}|Is6yd5o6b1ba,Ht;*8bIGjrBa3|\\\"\\\",2):f(\\\"\\\"{>=atj1b3eR:BpXaQ/0rt0ADcbqk=@0bW0A6v+fG:qHu2*7bD\\\"\\\",2):f(\\\"\\\"{Oabb*D5be+,FSAt3X5V=Z;R\\\"\\\",2):f(\\\"\\\"{B\\\"\\\",2):f(\\\"\\\"}<aD-G4*zb51b8>OL:/wb\\\"\\\",2):f(\\\"\\\"{qmbB>Lvub/-jA@a5o<aFDFo8bXa;0Wa0be,9bEa.,T9Q=O=R6AH?J.bdb7bhb\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"}BCYag,EaVaF2\\\"\\\",2):f(\\\"\\\"{8"));
$write("%s",("Wa/-4tVaubJ.jbN6c38|09L*W55oQtb|?F<a65vl?fDa:rI=3blhSag-FgK-kbUaN-ebXa:HB|a@iblG5o*xGDn21zPz+@\\\"\\\",2):f(\\\"\\\"{b:k*b..t0\\\"\\\",2):f(\\\"\\\"{b|u7/SwVa8b0|,bTaO+OaFqQxxIXaFai,8b3r/Ac1NaNHt5cb;:5omEvvIGwb1J1bjb*5hb/wcJQ*Z|,iKC\\\"\\\",2):f(\\\"\\\"{qY\\\"\\\",2):f(\\\"\\\"}IwPEhc0sAav:vbo|6blb4pHnr\\\"\\\",2):f(\\\"\\\"},0e0Eu6bKG9-\\\"\\\",2):f(\\\"\\\"{wvqSa8b4eSa>IYn<.x-ToQH/GFaubM\\\"\\\",2):f(\\\"\\\"{A?<..,,bQt:ppvhbU.*3q\\\"\\\",2):f(\\\"\\\"{5FAHH<oh>@pi+bFaEr2,i4/bRv01tbcbAwu;dx>agJ<aGal*+:BaBw.kkb;3X2Lq3\\\"\\\",2):f(\\\"\\\"}4GYgS2b*Sa\\\"\\\",2):f(\\\"\\\"}IPaQ3RvQ6Oazbyb*by?7bzbn7-6=B50kb/t1vfwQc-qB|n|l|4EakSaPtWaq;rgl4Va3b7Ieq\\\"\\\",2):f(\\\"\\\"}bt+:zDjg,U\\\"\\\",2):f(\\\"\\\"{avfbgb9;Dai61bgoBazy/byzfvYaebWaLE@aakB?r,ub|v.H0b\\\"\\\",2):f(\\\"\\\"}bA*Tan>m-s11kib\\\"\\\",2):f(\\\"\\\"{*ZyLpQ+k.bv;rq><uP/d4fb-bS2l+ToIH.bFaBfp,-*S2UoD\\\"\\\",2):"));
$write("%s",("f(\\\"\\\"{mb?vr2SaNjCt9bm-@aVab+mb.HUFA*4a?Hhn3F;FOau\\\"\\\",2):f(\\\"\\\"}sv9?5GZa?ak+GwD,hb\\\"\\\",2):f(\\\"\\\"}bp,<aq,zbvb1vjb4@SajbYaku,yXhiubbBa9?3zE*XoRaayMpHFLrIoHkT*jbkbYF@afw?aVa6+|bU5<ai*;q<mzbdb\\\"\\\",2):f(\\\"\\\"}zP/>qNFD3\\\"\\\",2):f(\\\"\\\"}bTo/be=@a7h23,pOa18\\\"\\\",2):f(\\\"\\\"{b:*s4cDE0@al=CaTasx*zqo</<a-GvbP6.12;Co=a5bFa9vmo*bzbavRaAa,i9bFa?a2\\\\\\\"\\\"),\\\\n(\\\\\\\"\\\"9I.PaT>R8>aXaMq2bdbn:|bawg-@a0b9rJ\\\"\\\",2):f(\\\"\\\"}5ob3Bam5BaXav4,bjbqwIgxv\\\"\\\",2):f(\\\"\\\"{b\\\"\\\",2):f(\\\"\\\"}-\\\"\\\",2):f(\\\"\\\"}4TafwEvOq@aav,bUC:/hb7q.bRvpttb4bC\\\"\\\",2):f(\\\"\\\"{lbav4bB?jny@i1R\\\"\\\",2):f(\\\"\\\"}+B,l/DNhWa*4hbUi,bjiZDF23b=3Yt7v*bPaauFaOaAat/n9Tal9j9ub,yk>cxpEkDDa;@hDXavbZxG4BC1bb6.3tbY,q2NaNozbPaXaay\\\"\\\",2):f(\\\"\\\"}b.bXaB9soA,wbC>RaTrA*>\\\"\\\",2):f(\\\"\\\"}mbFz8b\\\"\\\",2):f(\\\"\\\"{btbCavbLru7hbZaJoJdGaN@n8Ya5bWmWawbHyr@"));
$write("%s",("jdn|dbtbmw9bc66CJ9O=NaAtFazAd.\\\"\\\",2):f(\\\"\\\"{byboj8be4ovl7S,y:/-ICSaYa;A=aG/h>DrKC4pxb9t7bPaTaWaE,ecv45s3bab7pf=kvAu?a6+eof-92vf:\\\"\\\",2):f(\\\"\\\"}+|:\\\"\\\",2):f(\\\"\\\"}7vhb2bvbg\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"{bx|gjNj5wPuj1x><x\\\"\\\",2):f(\\\"\\\"}BnC<:x-suXa=zRzwbm+5oF.W5ld4Aoxbb<aQvKC8b31k+5;fbr-Wvq3|w>uzbs6Oa>@7bSz,\\\"\\\",2):f(\\\"\\\"}lov93bjbJ0xbab3:ttKrqtl9y:aberUaGtP>=an<ibib5b6t<aYa+yJ65<*b+p+uc60b0y8BYaZ:Rv|z|bT@Ua\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"}*<C*2b>aC*2xR8sji:IwUa+bN8Xw,b7r|b0bZak+ewqr6.aoABUa1o.,zbd77*9b6b:zdbBaUa@,hbUaj+@a:zD3Takbxbg7zb.\\\"\\\",2):f(\\\"\\\"}rg+b,qGax=A*e=RaD,-b<,Na>a2zU\\\"\\\",2):f(\\\"\\\"{8beb,y9b+pkbVtCwCA@,Puf1s<4lD54l\\\"\\\",2):f(\\\"\\\"{@zb0v/bHAfxR,5b9+t+AfR:BaC2UvZaw;qsCiaq9*+p</Ta5ojbH@q0zvy,\\\"\\\",2):f(\\\"\\\"{bY*hlq3jb5oyb5<d,+y8q1-m1E6-sbbKyD,fh.x8gUY2y-b?5d"));
$write("%s",("g8w.,B;eq@*,br,zb2<gxtbswcbuu.z+ber\\\"\\\",2):f(\\\"\\\"{bab|w.beb*1n>Jvib>hgb6/8-ck=ax-8g>uyb=0\\\"\\\",2):f(\\\"\\\"{bZbXa+b8b<a?aTt7\\\"\\\",2):f(\\\"\\\"{Vauv50x4|bMwubf?tbzb*?Wafycb:=ib/|jiB/l=@8.3P+DoWaXajb|u-bWaAaeb?5/b-ba4@a6b,\\\"\\\",2):f(\\\"\\\"}B6tv5btbWavbz+j9U|qozbTa|b?\\\"\\\",2):f(\\\"\\\"}UaW\\\"\\\",2):f(\\\"\\\"{Ya1lx@IbZ.v>Uaqk>atbzs7b,7Aawbtroyjij|3gM.oyl<;?+*tbZ7:7QaW\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"}m=ae<ovmb=?qkRa,7X|4;r\\\"\\\",2):f(\\\"\\\"}lbC=FaxbN*Fam6@-Eac-Wacb|bGzXlk.>a2?8b>vwbz;kbFaeuZ+mzazQxzdns<9CaZb*>\\\"\\\",2):f(\\\"\\\"}b0j-b.to>7bgbX\\\"\\\",2):f(\\\"\\\"{t?gw7\\\"\\\",2):f(\\\"\\\"{6w<tw,R:ixau5\\\"\\\",2):f(\\\"\\\"{<aQ1+x1-6b3vSal7OaT9\\\"\\\",2):f(\\\"\\\"}b|b7\\\"\\\",2):f(\\\"\\\"{7vxbW8e/TatbZhJom\\\"\\\",2):f(\\\"\\\"}Qa2=\\\"\\\",2):f(\\\"\\\"{ovbSzC0PaB6W67-cbT9gbGyjb;tibL;>uWvQao7L-jdlbcbs\\\"\\\",2):f(\\\"\\\"}av.vIsAaPaRanoAa9bL*f\\"));
$write("%s",("\"\\\",2):f(\\\"\\\"}SahuZqXtPuT\\\"\\\",2):f(\\\"\\\"}c:T7p<A\\\"\\\",2):f(\\\"\\\"}W0P9hb@a9b\\\"\\\",2):f(\\\"\\\"{bmbcb*pab.x\\\"\\\",2):f(\\\"\\\"}bmb>w/qxqqxl0j0,sabfyYaXaCp/be5=w55b5/blb\\\"\\\",2):f(\\\"\\\"}bQaaqCt0bD+rzytdx@aO4ZaXa4b0wcbxbttXlB;Xa2be03b@t6u\\\"\\\",2):f(\\\"\\\"}omslbjb+-fqxq|5fyo\\\"\\\",2):f(\\\"\\\"}gbb-h+fhubjiN/PajbW|Q+5otbJpzv=|\\\"\\\",2):f(\\\"\\\"{b.\\\"\\\",2):f(\\\"\\\"}7bZsWaf=p:gbkb+b4*ZtTo50U8GaO7Mw7buyK9Lu/8w9Q0Vpb0=aDv..t,m<7bp;X/ksMmn<Hwb<I+z8WaSaOr?a7blbJ./bp;|b9+|bRaVaTalsJ.\\\"\\\",2):f(\\\"\\\"{yksTa=aFqS1Iq6qo|SzTi9p1lY.F5s\\\"\\\",2):f(\\\"\\\"{|3a:WaTa@a>qqrf<r.Mrmb@-PaWa@aSaMmOaVop:5o3bwbsy2obrs9*bcblbTpvbBapxO,-4ub-6ab1x4bTikb1b<aabix5-OaSayb\\\"\\\",2):f(\\\"\\\"}b?a\\\"\\\",2):f(\\\"\\\"{b5b2b.b0bYa47hxfyat7\\\"\\\",2):f(\\\"\\\"{Aa0bO,3svomb0btr|b9bRabb|bQqUvkb8r0h47lbqrHtQam3ztdbhc0|lbmvab|bH-\\\"\\\",2):f(\\\"\\\"{b1hW5n8Q"));
$write("%s",("tH.fbCaXyhbQqoyGw\\\"\\\",2):f(\\\"\\\"{yyy5bitBzUa=iQt0+d9bvy:Ea1bZqP1Va=aQaY8a*i-Uawb\\\"\\\",2):f(\\\"\\\"}bOatb-0Rawu6bEj9bmvkbsp|bNpibJ6d38b+p02gb2*OaXa;zlbFib\\\"\\\",2):f(\\\"\\\"}-bZaNaMqjiAlPu>x\\\"\\\",2):f(\\\"\\\"}3*,U7Va?aOat\\\"\\\",2):f(\\\"\\\"}*bfwvb>,\\\"\\\",2):f(\\\"\\\"}sLsvbTaPa*wrgwbPasoHrBrpqGgtjW5gmb,hb5zibg\\\"\\\",2):f(\\\"\\\"{8b+exb@u<uL-\\\"\\\",2):f(\\\"\\\"{5E/dgOaybLnwbhb.qEuHy4ubbpp7+JoJu>\\\"\\\",2):f(\\\"\\\"}p+2bDaC1+b7bxuvbib=aybF2TpDaPaYamy=ic*4yE8|bmh=avrT3Jwp6gyxbRa-vOas/98FiNaO\\\"\\\",2):f(\\\"\\\"{5oBa6bUyS4ZyUa5bVa967bFizb1o>.7rJqTo/tFa4b=agbZa@qA,n|jbR*DaX|*byb1bSaPamblbVaVaOas+YaEa:4Gw8b4b0|tbab*|*qUak2o7m7uoFazpWm2xNj2xEa\\\"\\\",2):f(\\\"\\\"{bC7hqjnR7C5V.A5@70o>7Z-fbI5n2ewEq/-Ew1bDaEq7\\\"\\\",2):f(\\\"\\\"{aocb5bt5vbA-vbk0>aabkrh\\\"\\\",2):f(\\\"\\\"{gvv75b/bub1jE,Pq>qsrwb>aR6KtB|zb\\\"\\\",2):f(\\\"\\\"{bgb02abbb"));
$write("%s",("hb4bBaXlAaE6,bSaXy7b>\\\"\\\",2):f(\\\"\\\"}x35qV6Uaw2h\\\"\\\",2):f(\\\"\\\"{|bntN69fOa*b82FaMw-bL4p,ybhb,bUaab/6vySavbebebBaNa5b5u+4ab0bf\\\"\\\",2):f(\\\"\\\"}fb\\\"\\\",2):f(\\\"\\\"{6pz;kDan|>aFohhRaNzZ0\\\"\\\",2):f(\\\"\\\"{zkb5->axb+-6b4wB\\\"\\\",2):f(\\\"\\\"{4s7\\\"\\\",2):f(\\\"\\\"{|utb9-\\\"\\\",2):f(\\\"\\\"{|ib|s=a+cdb.bAaIwlbFw,dVaFaVa8rXaTaJn0wVattZalb\\\"\\\",2):f(\\\"\\\"}orodbXaab6|zb7sAaubBxyz+x=t;tVwcbGnAas\\\"\\\",2):f(\\\"\\\"{,,8x1lP\\\"\\\",2):f(\\\"\\\"}U.N\\\"\\\",2):f(\\\"\\\"}z32pUa-uibSayz.wtb@fAaxbxbcx8blbQaI,gbAa/bjbgbCaNaebVa9wsoW24s5bto5o5bib5pToEaybwbAflbwbys-b6r>aTa@\\\"\\\",2):f(\\\"\\\"}NpabWai45g6b4rybyb\\\"\\\",2):f(\\\"\\\"{szb=zNaJ08b.d0box4|vb7z\\\"\\\",2):f(\\\"\\\"{uab5pybWaPqAse+/bwbW|BtzsW0Xa=aJ-A-Oa@aDaAuOap3?2GaL/6bEaebPa5bso+\\\"\\\",2):f(\\\"\\\"}9ik0=u4b*b0b23mbbb?\\\"\\\",2):f(\\\"\\\"{,bkbZu6bDaeb2bebN0lb=t<m2b1b4r8bh\\\"\\\",2):f(\\\"\\\"{z"));
$write("%s",("bdxtb2b+bkbQaQa0b,d-bDcFt7b>aUaotb0\\\"\\\",2):f(\\\"\\\"}be+5u6b,+k,,b1orz<3eb1bGaTwvb7uc\\\"\\\",2):f(\\\"\\\"{SnSa*bD\\\"\\\",2):f(\\\"\\\"{2bZhdbldXacb.ks\\\"\\\",2):f(\\\"\\\"{Tuh1W.\\\"\\\",2):f(\\\"\\\"},e1soQa*rF2*zcbZ2CaQa8b6b-bkbScD\\\"\\\",2):f(\\\"\\\"{.k>aS-Zatbwbvb7bDaFgib0o4,ibNlSa<.db3bl|voSyVpWaw0w+fbvbGuTaUa0bGp\\\"\\\",2):f(\\\"\\\"{bib1bg-2bj/7bU+Na|b@aUa/*tbD\\\"\\\",2):f(\\\"\\\"{ybmwwbFn.bcof0fb9b*b0s,\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{qkbW1@q9wt+k.Hvczcq/b|b4b<,/bm|AaNa.tauYabbM.ewI|3bgbTaKyMrUyr\\\"\\\",2):f(\\\"\\\"}.th\\\"\\\",2):f(\\\"\\\"{Oa4b*1huCaabI1?ymb7bO,Y|3oA1ji?1TyvbFaib5o=0OaNa.wxbtb51@uA,/sov+bwbmbfk@akb4bYa@.EadbDa3\\\"\\\",2):f(\\\"\\\"}-*1\\\"\\\",2):f(\\\"\\\"{K0xbi,<a1y<afb=ahbYa2b<akbk,jnU.r\\\"\\\",2):f(\\\"\\\"{S.RuziX.2bYa7-5|abYp\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"{3bO0;m+bl0-hFaCwNp@ahbgwfbXadbbborXaeb-bab,iwbVazbb*ybeb"));
$write("%s",("+bYyzb=u5|+b*bnt2\\\"\\\",2):f(\\\"\\\"{e0:+.b:-h\\\"\\\",2):f(\\\"\\\"{4b@aeoJrtb3s>ar0.bM\\\"\\\",2):f(\\\"\\\"{K\\\"\\\",2):f(\\\"\\\"{=a4p|bcrYawbV,1b=ary*b/b+p2ov+t+BaFaX/9y|bi|Ya|b2bXoA/PaA/P/yvQa>aG/OaJ/F/>aD/\\\"\\\",2):f(\\\"\\\"{pT,5oSaT,ji8,>aZ,a-ho,b7bwbGazx-.lbmbebo.e/J.>a1hgbTy6.BaIoRag/\\\"\\\",2):f(\\\"\\\"{/J.l/f/d/8s|s4bvb0bRam.k.XwJ.Xwh/Uah/QaVa-.jsq\\\"\\\",2):f(\\\"\\\"}Eaksut\\\"\\\",2):f(\\\"\\\"{lxi|,:x+,O\\\"\\\",2):f(\\\"\\\"}t\\\"\\\",2):f(\\\"\\\"{M\\\"\\\",2):f(\\\"\\\"}S\\\"\\\",2):f(\\\"\\\"}7xFc1h=yOalbPayb1hRa?ahx\\\"\\\",2):f(\\\"\\\"}b\\\"\\\",2):f(\\\"\\\"{bDak.<aWa6-dbCaBa1hBa.b5.6.>aFy6b\\\"\\\",2):f(\\\"\\\"}mG-Dn@a1b@aJ\\\"\\\",2):f(\\\"\\\"}Ra-bYaVaj-Ra6-wb/bVaPa>aEaAaOa=a1h5->\\\"\\\",2):f(\\\"\\\"{mb=aEalbgbPla.TaSa@agbNaSalbRa.bg,xbgbEaPaq,Sa0hYa0bBa=aIqEaSaWamb@aRaS*OrCaSa6-@aWaOr7bjb.bYaOpXaZa.bRaabNaGq+p0babFadbJnayvbsvdb5yD\\\"\\\",2):f(\\\"\\\"{ZtD"));
$write("%s",("\\\"\\\",2):f(\\\"\\\"{ibebCa3xPaEy@a/bHdKqjtyb,bjt6b*bPn6bZagtDn/bRaT,5bRa\\\"\\\",2):f(\\\"\\\"{bOa4p>a/bZaDa+yo\\\"\\\",2):f(\\\"\\\"}8b9*ZaAaqkkvwbUagbf+UaNazbxhOa+bT*S+@a?aGa>|<|5o/bhbh+.bNa?ajig+Da-bPu2l\\\"\\\",2):f(\\\"\\\"{,n\\\"\\\",2):f(\\\"\\\"{fnQ\\\"\\\",2):f(\\\"\\\"}L\\\"\\\",2):f(\\\"\\\"}fb7bP+mbvbOaWat\\\"\\\",2):f(\\\"\\\"}mb>aFaKtQawrYa4bUalbSaNaabzbUa1bVa|b>a1bUa2|EaNa*v.bkrRa1bn\\\"\\\",2):f(\\\"\\\"}l\\\"\\\",2):f(\\\"\\\"}TqdbRa8bWamy-b+b2rzbt*BtkvSa:+?\\\"\\\",2):f(\\\"\\\"{QxDq4bhbCt?aYa*b*va*Y\\\"\\\",2):f(\\\"\\\"}W\\\"\\\",2):f(\\\"\\\"}To3blbQx,babmbgu>\\\"\\\",2):f(\\\"\\\"}Afibzb:kuudb=a\\\"\\\",2):f(\\\"\\\"}b/bXadgQaEa5o+blbkbNa3b;k5o0blb-bL*;r<a;pTaNaU*M*?a*b>aOa,bdbUy.vjbOa3bdbUaPafhCaFa*b-sZa-vYaDa6bbruk=teb7babwbOaUaDawbebzbZa@r\\\"\\\",2):f(\\\"\\\"}bZaYa\\\"\\\",2):f(\\\"\\\"{bkbEaR|Ta0bLwttwbm|wuFztbtb8bmdPv3\\\"\\\",2):f(\\\"\\\"}?zji;|Ao=a5oVohb+o=i0bRt"));
$write("%s",("AavfxbCa5b*b1wjns\\\"\\\",2):f(\\\"\\\"{dscn9xo\\\"\\\",2):f(\\\"\\\"{s\\\"\\\",2):f(\\\"\\\"{m\\\"\\\",2):f(\\\"\\\"{p\\\"\\\",2):f(\\\"\\\"{k\\\"\\\",2):f(\\\"\\\"{EiUaXa0b1h>aP\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"{z9b=aib6\\\"\\\",2):f(\\\"\\\"}abubCafb*bQaCa;w9wWaDaY|,bubww4btrBa;pOafbcbTrbvkb5\\\"\\\",2):f(\\\"\\\"{RaZa*xLr*b=aYaRaOa\\\"\\\",2):f(\\\"\\\"}rZambwbwj\\\"\\\",2):f(\\\"\\\"}bAabbHnubzb+bfbXhyb8b=akbgb+b8q?pab3bZa4e3bFa-bhb>aa\\\"\\\",2):f(\\\"\\\"{2w6v?vxq<aub+cvb.bQy>alwvwvb5oFaurdbebjbAaBaeb|bhbbbbbNaLv-t@z/bEaZaeb>avbrsXa?va|Oag\\\"\\\",2):f(\\\"\\\"{UpybvyogVa\\\"\\\",2):f(\\\"\\\"}bSaub5oRaub*qbbF2RvcbEazbeb3sqotbTaxbK\\\"\\\",2):f(\\\"\\\"{bbOagy0s\\\"\\\",2):f(\\\"\\\"}bPa1b7bBabb-bAa5odb6bPa0bdbzb5oCaWaUa?a;uVtCaGaMxgytb\\\"\\\",2):f(\\\"\\\"}bBa*bZa4pBa8bhsQa5ofbFa:zufjbPaSaFa\\\"\\\",2):f(\\\"\\\"}bubXaPuQul\\\"\\\",2):f(\\\"\\\"{Oucs;xasPufsbs=xlbtbPawbor/b.bSaAwvbPz9b,bhbNab"));
$write("%s",("b=wjbZaaoXa2tRaCa+bMn5bNa:pwbNaTozz,bgb>vub3bio4bDakbPavbybeg4x/r-o5byb=aNa0b@tsrDagt?afbibwbXaRaeqcbusebwbyy,bEw2b@t/y3b;u1bIwSacb:yut@gabTa>qPabbYatbybkbOa/bDa1hXaDa/bAambjqlbXazbkbAa.bDaOa2bef8bPxzbRa0bkvOaTa?a2gzbro3bCa5o2bAaGu=aOa2rbb4b-uGwTaebSa3b9bcb8bmb1b+bmbEambgbUpBaFqitZq*bOaabib.bau6s1bcb3b3buw3b?a1boq9bmxAaauJxUwQwVwZqNa4p3bBatbzuCaautbBaaujnPuSugplpmpxikpPuan8vPa2b8bjbct1oPa>tnvkbmbjuhc0otx6b,bVvdbDr*bRaBa5b8b7b4b:q@t9b\\\"\\\",2):f(\\\"\\\"}b3bYacb/bOaubgbYtCt\\\"\\\",2):f(\\\"\\\"}b;r5ows-bji\\\"\\\",2):f(\\\"\\\"}t2bFs-b>vabufZaXuAa4bXambAa|bgb3bebNadb-bkvxq@abbubUa|bCa;tAaVa*b2bUaCa,b8bibAq<sGujb8vkbBaYahoMo5o1bbb+bgbqwcbXaEvcbCaji.o3r0qTaFa0bNaibRrib>a5ouk6bdb5bZa|rgvkbeb9btbjbab7b>rPakb/bevnowbEatbNaBams\\\"\\\",2):f(\\\"\\\"{b?a4bLtmbNp7bXaQakbab3qcb.bWaYa,b*bTabbcb"));
$write("%s",("Oaavtb\\\"\\\",2):f(\\\"\\\"{b/bcb6bkvgb5bOaCa=a=a2bTaab4bmbBaPc4q2q/bUacb9b|bYaQa\\\"\\\",2):f(\\\"\\\"}bIgbb@qCaPuYrNuZr4aes0lWrgbhbtreb<stbbbib2bjbdbcb+bbbxb0b\\\"\\\",2):f(\\\"\\\"{bubdb@q>srsdb,b+b4bgjEafg6bfbmb5o4r4bWaIn4bZa=a@aBaxb8bOa+pzbAaQadbwb,b,tbo0beb\\\"\\\",2):f(\\\"\\\"}bEaauubAa>aYs-dgbmb3b<aHtZa,tOacb0bcb=aUaubyb.bEa=awb7bdbVaco7pgb\\\"\\\",2):f(\\\"\\\"{bAatbbq7btbdb*bmbFaSaSa|bkb5o9bvb,bRa7bNaValbHr5o\\\"\\\",2):f(\\\"\\\"}bYaqk*b\\\"\\\",2):f(\\\"\\\"}bcryb?a3bTacbUp>pUaib,bebTaDjRa5b.bxbtrrqNa\\\"\\\",2):f(\\\"\\\"}bVatbfbwbSaXhib\\\"\\\",2):f(\\\"\\\"}bTatp8b,bFaogCaOaxbDa.blbbb6r5owrur4b+bTa*sosmsfqWazbbb7b0b,bWaCaebtb|bUaxbTa\\\"\\\",2):f(\\\"\\\"{bUaybZazbjbRahbTaub5r\\\"\\\",2):f(\\\"\\\"{bYalb9b.b?aeb@qubQa\\\"\\\",2):f(\\\"\\\"{b.bUaVa5bhbjnxiipXrjpnphpjnjnLibpQawjvbPpxbDjVaSaTaBacbmbmbXafbhb0b0b5o\\\"\\\",2):f(\\\"\\\"{bXa-b@aV"));
$write("%s",("i0bco@a-bfb|b6bjb,b-bmbjbcb@qYaub*j9bPa\\\"\\\",2):f(\\\"\\\"{bTa1bFa.b=aerFaQa1bfbOa8bUaQaSc,b:qUqlb7b5bkb0b8bjoebOa1bXa5q\\\"\\\",2):f(\\\"\\\"}b\\\"\\\",2):f(\\\"\\\"}b2q;q9q7qAa7bcbFa|b7b-bFa>a+bjbUaFoWakb9bVa\\\"\\\",2):f(\\\"\\\"{bRazbNadcub\\\"\\\",2):f(\\\"\\\"}b1bdb8b.bTaQambabebQa|blqjq>aNavb5b@aFa+bApFaNpLpvb1o-b5bDa1bub|bVadbOn\\\"\\\",2):f(\\\"\\\"{b@ogb4bjbNaMhkbRavbdbublbvblb\\\"\\\",2):f(\\\"\\\"{bebmbibTadbTa0glbabcbYaabYojbJo?ecbhbGoDazbEaEakbbbfbZajb-bEaabjbhblbYaZaeoDaDaCa*b,p+dXabb\\\"\\\",2):f(\\\"\\\"}b7g5oNa,bvbJo=a,bZahbDaxbcb?azidpep,lcp,lfpinzimnnnzilnjn9f-hjb>aebibOa0bibvbZafbAa5b3b\\\"\\\",2):f(\\\"\\\"{bcbwbabDaFa1b,b5bebegkbdbkdab9bwb*bCa7b|bDaGa/ogbvbNa1bjiqb7b<a>adbAalb,bYavowouoso7b/bYagbibjbDavbvbPaEa+dFacbgb.b-beblbzb,bNa7bvbCaEahb<aCabb*bohQaub*bWaQagbSa,bEa7b6bAaEaLl6nyn>mommmrnXfAmum0n;a"));
$write("%s",("Tmvm?atmTm@m>l*n-bLl7mCa=lQmwbicTm?llmunEaWlAmnm=l\\\"\\\",2):f(\\\"\\\"{mimgmjn4l4ldn4agn9axien,lbn/lzi3l/b\\\"\\\",2):f(\\\"\\\"{f-a:hub?h8a8mEm|mJm<l9aEaOaAm?m0m1i:a-bAm=aAa-a1m+mCaWlamzm@a<a-b|e4m*mOlkmZlQlOlMlrm\\\"\\\",2):f(\\\"\\\"}m:aCa|ewm>aAalmVlQl9a:lRlAa:kHl|ejmwlLlYlBa-aNlGlEl*bvbtb/b-a+bId@lSlAlJl@aHlLlSe|eFlKl?aAa=l\\\"\\\",2):f(\\\"\\\"{b;lBl@lFa>l<l:lHa8l9a|e9lxb8a+e-a1beg8aXftl8arb|eidwi1l1l-l3aKixi+l-fyimlNhFf6b-a+czbxbubHaqb6aqbDiEiCi5aqb@g-a,bAfzb.bKfnbxb|ijiZgXg\\\"\\\",2):f(\\\"\\\"{gag\\\"\\\",2):f(\\\"\\\"}h6i?kvh=ktcBa3a;dLfak@k3kVjBa?a3aOhIgCiwbJa7iChYj*hWjDa?a>aJi6e:hrbbkZjhk4jCaJi2b3bFiUfxj8f1iCj?a3jKa\\\"\\\",2):f(\\\"\\\"{b;a3gwbccIa3b1b,j,b|b0avh7hvhPiNiLi@aJiyb3bSj?a8j4i5h5jBaKiMf0i\\\"\\\",2):f(\\\"\\\"{g\\\"\\\",2):f(\\\"\\\"{gsbubwbji-aCjAj:a;b>j1b0b-b3aAa3a7b-aji.a:b:b,b7hVhOiliMi@a3a:hwb+"));
$write("%s",("b-aPctj/b8b1bPcxb;aUf-b:fZapg|b.b5b-alj=i3bWfvb|bIgFipgfg3bgf;a<b:b3b-a8bIg,bxb2b2btb;a7h*h5iPa3i3a>a3a5anb-aDi/b3b4b.bHa8byb2b2gtbWfxb5b+bYg7h5hkiXhVh;d+cKfHa,i,iFaGaii|fld4a.gvi/auh4a-afgdgMaFa=aVh-bXhChBhGa+bJdQh9a/b5a|fCc8g-bPaBaobChHfMa9aMaIa5axb3b.b4b0bxbzb-btbeg7hkg5hGaMbHg2bzb;azbLfccJaoh?auh*hCdYaOaVafbVaibNa=avhvh?a;aSgVaNaUa.guhkgvbpbEa*c7b?aCa>aDa>anbJdubSczbPfIcQgyfwfuf2bsfNd3bHa?e-a-fZf:aIa+c9f:avbldub4bcb-b3ggc0gHaebdbJaGagfef8a1bxbwbtbxbUaac|b3bdgfb/akgzgtbxcRf?a1akg-a6a5bhg>azd:a,cNahgwb.b;b>aagob,c:a-a.b\\\"\\\",2):f(\\\"\\\"{bvbxb5a1aob,fCe2b-a:b1dtbHa6a/c2b/a,fPcFf/b:b6aKa6e1b4eIa8btb1b1bNaGatb5a+ctb,b-a\\\"\\\",2):f(\\\"\\\"{fyb3dMd-aDdBd@dmf/aob5a.d,d*d-b4b7eSc;axb+b.bbcZb0cbfJasdHa/aed+e0cGb/d,btb-b4aWbudpcgdLc=chchd6areOapc0cNb/a;bje/eGaHb5dedOb.a"));
$write("%s",("8aNd8aLdLa=a>aIaOaJapb6a+e5azb+cdcfbhc;aOaFdYd6aHaCa@aIaQd8aHa=a.cIbCbMd\\\"\\\",2):f(\\\"\\\"{cycvcocRapcXbocTa;b;bpbgbYdJaGbRanbQaJagbnbcb>dqc5dpbebnbOa8a0c4aJaTa5a+btb5bxbJaQa,c*cRa5a1bzc6aedMa0c3bldjd;aeded8ard5a6a5aedxb/btbvb2bxb,c1b4b3bxb1b0cocPa8aNapcMagdUc3b|b+b/b2b4arcFbnc4a=a?axbtc4aSbJcPbKckcic+bZb3b-bzcXbqcFb5aMa/ancvc+b+b|byb4a9cVbNa5aRb7cFbnbFbMapb2c.aMaFb.a4a5aJaOa-a-b|b-aeb5\\\\\\\"\\\"),\\\\n(\\\\\\\"\\\"aicybHa<b/akc>a>aXb6aOb/a8a6a/apb4a1b.b3bvb4b1b3b2b-b.bvb4anb/aJaPa5a8a4a6apbEb5a5aBb,b9a4apbpbnb8anb4aGa=a:bJacb!\\\"\\\",2):f(\\\"\\\"})23(f\\\"\\\",2):f(\\\"\\\"{#~[2xha=s,y=z,13&X3^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):"));
$write("%s",("f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'yay,]99999[gnirtS wen=][c n3aea\\\"\\\",2):f(\\\"\\\"{)v]y3b&a(niam diov citats cilbup\\\"\\\",2):f(\\\"\\\"{RQ ssalcz4rfa cdlnl3c/a;maertStnirP/oi/avajL tuo/metsyS/gnal/avajm4bdateg@3doa2 kcats timil.v3dga]; V);Q4aC3ecaL[b5aX4hha dohtem?3e;4nga repus&3ecaRQ@3cgassalc.<5joa(=:s;0=:c=:i;)|4ajaerudecorp/3fqa(tnirp.biL.oken\\\"\\\",2):f(\\\"\\\"{.3bianoitcnufR6\\\"\\\",2):f(\\\"\\\"{sa(rtStup=niam^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^32^[2fha\\\"\\\",2):f(\\\"\\\"})1(f\\\"\\\",2):f(\\\"\\\"{#v3mja51(f\\\"\\\",2"));
$write("%s",("):f(\\\"\\\"{#,4353(ga13(f\\\"\\\",2):f(\\\"\\\"{#j4[j4boa(etirw.z;)tuo.N8aba(67b~auptuOPIZG.piz.litu.avaj wen=zG4Zka30341(f\\\"\\\",2):f(\\\"\\\"{#tm4[m4c5aR0Z0Z/512152353/2/2166263=4/3141726??:1518191:1/@4[@4cda*6 Q5[p4dea1312^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'5[w8[$5ofa41310r4[r4c7=[B>[j4[^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'6pma(amirpmi oicy4[(5[j4hma++]371[]591[?6[?6cpani;RQ omtirogla\\\"\\\",2):f(\\\"\\\"{4["));
$write("%s",("\\\"\\\",2):f(\\\"\\\"{4cCa;t:\\\"\\\",2):f(\\\"\\\"}%%%%\\\"\\\",2):f(\\\"\\\"}fi\\\"\\\",2):f(\\\"\\\"}*-84\\\"\\\",2):f(\\\"\\\"})48361(f\\\"\\\",2):f(\\\"\\\"{#]i[\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"}+17\\\"\\\",2):f(\\\"\\\"{<84.;i:-i602\\\"\\\",2):f(\\\"\\\"{;i:911\\\"\\\",2):f(\\\"\\\"{;j:632*7[ra116(f\\\"\\\",2):f(\\\"\\\"{#(tnirP.tmfIIcfacnuf;&4[&4bdatmfn4[n4cgaropmi;ILagagakcap~4Zea5102T6dbapD6[r4cba-l4[l4bpatnirp tesn\\\"\\\",2):f(\\\"\\\"})420aEaka etalpmet.r8[ma99(f\\\"\\\",2):f(\\\"\\\"{#(ntnire8[ia974(f\\\"\\\",2):f(\\\"\\\"{#fp4[ga^64^\\\"\\\",2):f(\\\"\\\"})32u9awa,s(llAetirW;)(resUtxeTOPada=:s%8[ba9#8eo4[ia9(f\\\"\\\",2):f(\\\"\\\"{#S Cm4[-Eaca&(y5[ga9(f\\\"\\\",2):f(\\\"\\\"{# .6[.6[.6oiaRQ margo&5[t4cjaS D : ; R-5[6L[j4[j4o%6[k4aqa. EPYT B C : ; Az4[56[j4[j4nka)*,*(ETIRW/6[J7chaA B : ;s4[s4aba [2cr4[*5dia: ^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\""));
$write("%s",("\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"' ohce3B[EYaeastupLRcdatniy4/ca0153.ea%%%%m4[m4[53ipaparwyyon noitpoz4023[230ca(nRO.%a7(f\\\"\\\",2):f(\\\"\\\"{#(etirwf:oin\\\"\\\",2):f(\\\"\\\"})4(f\\\"\\\",2):f(\\\"\\\"{#>-)_(niamp3cvP)ka(f\\\"\\\",2):f(\\\"\\\"{# cnirp,L)k;eja.OI[p]^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):"));
$write("%s",("f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'[(3rba@2Wa6;alaM dohtem06x*3c|5aU;cpadiov;oidts.dts 6Yab4kkaenil-etirwb5dva(,^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'s%^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'(gol.elosnoc;)^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):"));
$write("%s",("f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'73g\\\"\\\",2):f(\\\"\\\"}a^129^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"' nioj.)1+n(yarrA>-)n(=fI3cwa^31^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",2):f(\\\"\\\"}54,1\\\"\\\",2):f(\\\"\\\"{.^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"# qes-er()|3cH3bba^31^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"p3lg3fw3hla1% ecalper.j4dea^128^jAc/arts(# pam(]YALPSID^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\""));
$write("%s",("\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\".NOISIVID ERUDECORPA3cma.RQ .DI-MARGv3g53d|bNOITACIFITNEDI^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"[tac-yzal(s[qesod(^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"))System.Console.Write($^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"Put caffeine \\\"\\\",2):f(\\\"\\\"{(int)c\\\"\\\",2):f(\\\"\\\"} into the mixing bowl.^64^n^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");M3pva^"));
$write("%s",("63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"Liquify contents ofE3oeaPour^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'3w^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'4e\\\"\\\",2):f(\\\"\\\"{abaking dish.^64^n^64^nServes 164cma\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}^31^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");\\\"\\\",2):f(\\\"\\\"}/****/e3a^15^\\\"\\"));
$write("%s",("\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"),s[999999],*q=s;int main()\\\"\\\",2):f(\\\"\\\"{int n,m;for(;*p;)\\\"\\\",2):f(\\\"\\\"{n=(*p-5)%92+(p[1]-5)%92*87;p+=2;if(n>3999)for(m=(*p++-5)%92+6;m--;q++)*q=q[4000-n];else for(;n--;)*q++=*p++;\\\"\\\",2):f(\\\"\\\"}puts(s);return 0;\\\"\\\",2):f(\\\"\\\"}^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"))\\\"\\\",2):f(\\\"\\\"{s+=^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"00g,^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";for(m=1;m<256;m*=2)s+=^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"00g,4,:^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\""));
$write("%s",("\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"+(c/m%2>0?^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"4+^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\":^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")+^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\",^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";f(s);s=^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"4,:,^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";\\\"\\\",2):f(\\\"\\\"}f(s+s);for(c:Base64"));
$write("%s",(".getDecoder().decode(^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"kaAREREX/I0ALn3n5ef6l/Pz8+fnz58/BOf5/7/hEX/OZzM5mCX/OczmZzBPn5+X/OczMznBL/nM5mZzBPu++fPPOc5zngnnOZzOZgnBMGAW7A==^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"))\\\"\\\",2):f(\\\"\\\"{c=c<0?256+c:c;for(i=0;i++<3;c/=8)f(c%8);f(^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"8*+8*+,^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");\\\"\\\",2):f(\\\"\\\"}f(^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"@^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");^1^\\\"\\\",4):f(\\\"\\\"'|sed -e^1^\\\"\\\",4"));
$write("%s",("):f(\\\"\\\"'s/^16^/^32^/g^1^\\\"\\\",4):f(\\\"\\\"' -e^1^\\\"\\\",4):f(\\\"\\\"'s/^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"/^16^q/g^1^\\\"\\\",4):f(\\\"\\\"' -e^1^\\\"\\\",4):f(\\\"\\\"'s/.*/print ^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^8^nquit/^1^\\\"\\\",4):f(\\\"\\\"'^3^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")\\\"\\\",2):f(\\\"\\\"}^1^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")\\\"\\\",4):f(\\\"\\\"');\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\").split(\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\","));
$write("%s",("9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",64):f(\\\"\\\"^\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");for(int i=1;i<a.length;a[0]+=a[i+1],i+=2)\\\"\\\",2):f(\\\"\\\"{a[0]+=\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",89):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\".repeat(Integer.parseInt(a[i]));\\\"\\\",2):f(\\\"\\\"}System.out.print(a[0]);\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";FORiTO UPBtDO INTn:=ABSt[i];print(REPR(50+n%64)+c+REPR(50+n%8MOD8)+c+REPR(50+nMOD8)+b+\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"J\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"+a)OD\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\""));
$write("%s",("\\\\\\\"\\\"while(!=(S:length)0)\\\"\\\",2):f(\\\"\\\"{\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans c(S:read)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"D(c:to-integer)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 35 39\\\"\\\",2):f(\\\"\\\"}\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 24 149\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"interp:library\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"afnix-sio\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans o(afnix:sio:OutputTerm)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"o:write B\\\"\\\",9):f(\\\""));
$write("%s",("\\\"\\\\\\\"\\\");end;\\\"\\\",1):f(\\\"\\\"\\\\\\\"\\\")\\\"\\\",1):f(\\\"\\\"nsys.exit 0'}\\\\\\\"\\\")\\\"\\\",0)]]></xsl:template></xsl:stylesheet>\\\":s.WriteByte(Asc(c)):Next:End Sub:End Module\")\nput=s\nprint\nqa!"));
end endmodule