module QR;initial begin $write("%s",("let s=(\"Module QR:Sub Main():Dim s,n,i,c As Object:n=Chr(10):For Each c in\\\"<?xml version='1.0'?><?xml-stylesheet type='text/xsl'href='QR.xslt'?><xsl:stylesheet version='1.0' xmlns:xsl='http://www.w3.org/1999/XSL/Transform'><xsl:output method='text'/><xsl:template match='/'><![CDATA[sub f(s$,n)print(s$);:for i=1to n print(\\\"\\\"\\\\\\\\\\\"\\\");:next:end sub:f(\\\"\\\"write,format=\\\\\\\"\\\"%s%s%s%s%s\\\\\\\"\\\",\\\\n(\\\\\\\"\\\"\\\"\\\",2):f(\\\"\\\"write{-}{txt}{echo -E $'(\\\"\\\",1):f(\\\"\\\"\\\\\\\"\\\"with Ada.Text_Io;procedure qr is begin Ada.Text_Io.Put(\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"interp:library\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"afnix-sio\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans O(n)\\\"\\\",2):f(\\\"\\\"{trans o(afnix:sio:OutputTe"));
$write("%s",("rm)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"o:write(Byte(+ 128 n))\\\"\\\",2):f(\\\"\\\"}\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans f(v n)\\\"\\\",2):f(\\\"\\\"{\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"O(+(/ n 64)107)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"O(n:mod 64)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"O v\\\"\\\",2):f(\\\"\\\"}\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans D(n)\\\"\\\",2):f(\\\"\\\"{if(< n 4)\\\"\\\",2):f(\\\"\\\"{f(+(* 6 n)9)48\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{if(n:odd-p)\\\"\\\",2):f(\\\"\\\"{D(- n 3)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 27 48\\\"\\\",9):f"));
$write("%s",("(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 36 11\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{D(/ n 2)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 21 48\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 48 20\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans S\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"STRINGz:=REPR226+REPR153,a:=z+REPR166,b:=a+\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"2\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"+z+REPR160,c:=b+\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"8\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"+z+REPR165,t:=\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"#include<iostream>\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\""));
$write("%s",("\\\"\\\\\\\"\\\"+REPR(10)+\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"int\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"+REPR(32)+\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"main()\\\"\\\",2):f(\\\"\\\"{puts(\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"class QR\\\"\\\",2):f(\\\"\\\"{public static void main(String[]a)\\\"\\\",2):f(\\\"\\\"{a=(\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"write(\\\"\\\",4):f(\\\"\\\"'implement main0()=print(^1^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"BEGIN\\\"\\\",2):f(\\\"\\\"{print(^3^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"echo ^1^\\\"\\\",4):f(\\\"\\\"'f(s)\\\"\\\",2):f(\\\"\\\"{System.out.print(s);\\\"\\\",2):f(\\\"\\\"}s=^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\"));
$write("%s",("\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"389**6+44*6+00p45*,^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";for(c:(^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"#include<stdio.h>^8^nchar*p=(^15^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"Ra#include<iostream>^16^nint main()\\\"\\\",2):f(\\\"\\\"{std::cout<<(^31^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"class Program\\\"\\\",2):f(\\\"\\\"{public static void M83abbSystem.Console.Write(^63^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"Quine Relay Coffee.^64^n^64^nIngredients.^64^n^63^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9"));
$write("%s",("):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");for(int i=9;i++<126;)[3pva$^63^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",2):f(\\\"\\\"{i\\\"\\\",2):f(\\\"\\\"} g caffeine \\\"\\\",2):f(\\\"\\\"{i\\\"\\\",2):f(\\\"\\\"}I3b54rja^64^nMethodv4f#aeach(char c in(^63^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")))^127^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")^127^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^32^[2al3dp3c[2cs3c,3l[2k@3kqa^31^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")s rts(ecalper.h3eja^127^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f"));
$write("%s",("(\\\"\\\"\\\\\\\"\\\"     53c4a SUTATS(egassem^127^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"rts(nltnirp(])]^127^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\".NUR POTSu4cba.C3dh3dX3bba[65bX4df5lp3lna\\\"\\\",2):f(\\\"\\\"})1(f\\\"\\\",2):f(\\\"\\\"{#\\\"\\\",2):f(\\\"\\\"};)06xt3dba;+3noa3(f\\\"\\\",2):f(\\\"\\\"{#qp]\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"};)0,#3rv3rR3sv3mba723284-fa(f;)1q5.ba.>4[ga#(f;)3P6[=43ba7=4.<4[<4[<4[v3gJ=d=4[73++>u?4[73xda,43?4[?43ma^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"' D ; EYB RCo8[.6[?4;ba5qB/daDNE&6[&6[&6[8Emca AL9"));
$write("%s",("[)6[)6[v3oeaPOTS^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'6[^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'6[^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'6[M9pL9[(6[(6[v3moaRQ margorp dne16[16[16[v3lbaST9[&6[&6[JQ[~6[?4Nb"));
$write("%s",("a4~6[~6[~6[~6>ba&g=[$6[$6[.@neaPOOL|N[,6[4@[>Xp>4[#6[#6[#6[#6[#6[#6\\\"\\\",2):f(\\\"\\\"}da&,)l=[^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'6[^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'6[eUnga. TNUO9@[,6[,6[83nearahc1G[)6[)6[R9ogaB OD 0hU[-6[-6[%No33)$6[$6[%NBca)Av=[&6[?4<ba31XXk4dba0j4[fa#(f;)cT1YS[=8[*?[v3nqaEUNITNOC      0136[36[36[-FnV9[&6[&6[&FobC[^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):"));
$write("%s",("f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'6[^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'6[G@sba.)6[)6[)6[@4mja1=I 01 OD-6[-6[-6[C@neaA PU*6[*6[*6[v3:~6[~6[mTBxa;TIUQ;)s(maertSesolC;))T4[96[?4:ca11Y9/fatiuqnq41ca82p;[57[57[?4jda932A4.172ca65m4/i<[27[gC<ba9D?/maetalpmetdne.>72da215>7[>7[>7[?4kca007?/ca\\\"\\\",2):f(\\\"\\\"};^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121"));
$write("%s",("):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'6[^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'6[qD<ca66ZBWl4dba0j4[ga#(f;)4SA1batX6[=8[?4:da814>HX>8[cCkda283m4[x5[57gca0957/%a315133A71/129@31916G21661421553/:9[\\\"\\\",2):f(\\\"\\\"{;[?4:da378\\\"\\\",2):f(\\\"\\\"{;[b9[\\\"\\\",2):f(\\\"\\\"{;[x5[57wba5Q?0ra%%%%\\\"\\\",2):f(\\\"\\\"}*+1%%%%811 -;62ba5;D0;6[T8[x5[j4Fda21057/haj:+1 j@w?[W@[?4:da497W@[D8[b;[x5[b;wca3557/baww9[W:[?4:da082ZB[>8[W:[x5[j4vda6402?XV:[V:[?4nca67V:[=8[V:[x5[j4vda955l4.baWv9[V:[LX;ca52=8[=8[V:[x5[57ww9/ba\\\"\\\",2):f(\\\"\\\"{u9[U:[?4:da937<8[<8["));
$write("%s",("4Xiba4x5/wa)(esolc.z;)][etyb sa)^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'s7[S8[?4:kT0#6[#6[#6[#6[#6[7GM6G[;?[6G[x5[x5[x5[x5[x5[x5[x5[x5[x5[x5[m4[x5[x5[x5[x5[x5[x5[x5[x5[x5[x5[x5[x5[m4[x5[j4dda888iT[iT[iT[-W[#6[#6[#6Rba,%6[%6[%6[E9[#6[#6[#6~ba!m41ba6m4/ca~~37[37[37[S:[#6[#6[#6~ea(rt.(6[(6[(6[H9[#6[#6[#6~ba)BA[v3cda\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"};p4[SBfdadnes4[s4gra~~~~PUEVIGESAELPnr3ala~~1,TUODAERw3a:4[:4i$a(etirw;\\\"\\\",2):f(\\\"\\\"};u=:c;))652%%%%)u-c((||54[54ida#-<u4[u4ida||i15[15lhaBUS1,ODz4[^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\""));
$write("%s",("\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'8pka)3/4%%%%i(g:c4;[04jr;[r;wPa2=:/t;2%%%%t+2*u=:u\\\"\\\",2):f(\\\"\\\"{od7 ot0 yreve;i-=:u;1=:+i\\\"\\\",2):f(\\\"\\\"{od))1(evom(dro=:t elihw?s;)s*z9[L;ny9[y9uz4[z4i0Adladohtem dne.s3dganrutern3dCaV);gnirtS/gnal/avajL(nltnirp/maertStnirP/oi/avaj lautrivekovniJ3d25[25i[2cib\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"};0=q;)]q[c=z(tnirp.tuo.metsyS;)0(tArahc.y+z=]++n[c;y:]q[c?n<q=y\\\"\\\",2):f(\\\"\\\"{)0>2%%%%++i(fi;48%%%%)31-)i>3c&as(+87*q=q\\\"\\\",2):f(\\\"\\\"{);60212<i;(rof;n)rahc(+O5[O5q[2k.4[.4%oa=]n[c);621<n++z6aqa0=q,0=n,0=i tni;R4[R4%mc6ahi4asdRbQeelxfvfXk?f<bedRb\\\"\\\",2):f(\\\"\\\"{ke6;agb-a|dzdxd?fGb8aqeRdYd5aH96i;agb-epb>aqe"));
$write("%s",("RdHa>aJaRaAdteFbae:b6aOa5aacsgAzG89adL4aLa7a;a4a<a>hemkdxd;aNa?c6a|eebHaFaIaebzeJaeb9a/a6a2dQbUe-f2a-f9adL5d6cRbC3gdd-f/aof0f?fSg5a+h5e-,2e6aRa;dNaygQY1b6h;aTapc4aLcEehiof6amc6a-f;f<lsbdhrSDfybxcxc>aGaUeAa2a6ajg7a6a@ahg:a?aMbKaKa6a?e:aC,2aigGfMbIfUh>a:b1angcmBf\\\"\\\",2):f(\\\"\\\"{bHa4atc3bU,38k|+bsjk|\\\"\\\",2):f(\\\"\\\"}bJaMa\\\"\\\",2):f(\\\"\\\"}bJatLEc-bJaJaUa-bJaMdJa8bO7;a8bB-Ka8bB-8bTasj\\\"\\\",2):f(\\\"\\\"}bDPSaSa6+9bKaaINa?aTa8bwzB-8b6+<TJaLaJa8bwz6+n4cma8b6+4b6+:bk|,4cga\\\"\\\",2):f(\\\"\\\"}bJaHa\\\"\\\",2):f(\\\"\\\"{3aca<Tk3a)aFdL=;aaIUa:aUa:aO7ei@f>fDl4a/Qsbsb2be3^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\"));
$write("%s",("\"\\\"'maeiDa-a|b\\\"\\\",2):f(\\\"\\\"{*-aD6asaoHUe>awjhgKaKaigGf&6cgaHf@jRf*6esasbdh*b-a/bxcHa|f;1e3c-a\\\"\\\",2):f(\\\"\\\"}bhgXghgcg1ang\\\"\\\",2):f(\\\"\\\"{bHa;1?f-e:a:a\\\"\\\",2):f(\\\"\\\"}bHa?ahgJa\\\"\\\",2):f(\\\"\\\"}b=<1ba0<<.ec5aAdte@a1angsi;1xcpb7anb2b:bhg2f/j@dCf6aOjxcHaSfQfOfWj-aBfsigi?f-fng@f|f;1zeAggiHaMj;a/a3h<bmhFh<apb/a3hFhnbbM7b:bhg/awh:fnglgFaoi|b1aUh3b:bhg\\\"\\\",2):f(\\\"\\\"{hHa;1HaUepiCe|bxc3b0a:bhgIa|bzeJa|bc5auaQbgi<b=a-a;m*c3bxdUem3aea|b9ai3eta2bMa7apbuNXgVgTgRg9m3hCaAdI.Pcgfvfxbydzb7auN+k\\\"\\\",2):f(\\\"\\\"}kMa;m*cEc,dJa>a2a:b6ahjzkMa;m|b+i+cKh6a13g[a|b+i@JhVyg/a3h=aYhRaR-CdR-kbX+axYh2kEh7b5aMj?fwbkjUe2b5azgGi4b-bhcYrSjSjLu0c/bxd,h*hWi<@aea6a2bf@escvBfX6a|n2a5a,l+Jjg4hSk=vyjEhChinHa1dmd:h?f2k<kHa:e2k<k-l<b3bxd6a+h6k>hzljbThThvftfQY;aFicc35pbubldic+d,bnbWfcjajEc,d?a|jIkchGkvj"));
$write("%s",("<b<b<b5j:b+j<b<b,c:j7j7b-b:jKDAg3bDdvk<i9a7bwg-a2X,b,c:j=a9\\\\\\\"\\\"),\\\\n(\\\\\\\"\\\"a7bnuq3e13eca2j13ecaykA3c/3ggaJb7bKfQ3g\\\"\\\",2):f(\\\"\\\"{a1,Fj9a3?xb-a2Xf-kkXi5k,c:ji3a=a-aJdZVNg,c:jsb?fUjRk;k;i3jCa;i6aUjRkRjvj6aJk1kIjQktk<bzeVDceaHajgK5cca-k53c1a;k9k3a6a<bThKi*J2b2a2a2HOjLksiwbkj?f@a>anc:eOAa=aub\\\"\\\",2):f(\\\"\\\"{h5aDf=anbOjybok5a,bJa6a7b5aCgwbkjHa:e-b9a9b9aZjOjfg>am3a\\\"\\\",2):f(\\\"\\\"{a@a@aOjfg@a>a:a|b9a0b9a@a>aUCa?a>e|b>g9bJa0bOjfg-b9aZj9aCaAaJa9bOjnbJa6a|b5a,b?f:e-b+kZu-aW;a&aLu.JyNei2Hfg8bAd6h-a2H*b-.-a2Hfg7s3h5a2HKc-iA\\\"\\\",2):f(\\\"\\\"{xd6a-b9a8b9a7bJcJayb|m>aTh>aJa*c@dxc?bF0o3a5a-b;lteUe@a>a<a2bKdX\\\"\\\",2):f(\\\"\\\"{vb:atcJaub5aEcxbvb?a,b4b-bDgS7akaRjEk3amd:h17goaPkNkpb;awbkjplo5atb.JaZ,JYYJdHdrlyn<n5lYl,n*nwnk./n1EhbkoRaub4p8udb@S/w9xxRV+gsV+\\\"\\\",2):f(\\\"\\\"}bT,yvYsWym"));
$write("%s",("RSaJ9iR2+l\\\"\\\",2):f(\\\"\\\"}GGHncRRaTaX>HnU.WQmrG5p4a(day?tVn5bB\\\"\\\",2):f(\\\"\\\"{gb\\\"\\\",2):f(\\\"\\\"}w>4VBDa>4DavbhbN=Daf\\\"\\\",2):f(\\\"\\\"}/0I7kdWzvowp,o\\\"\\\",2):f(\\\"\\\"}s61GolPdF@a6pMGtbNpnPz2ZN9QI+sp2b=atbb+AvzD.1tLuwF|6/eb/b=aEalbc0gy/7;<<B,d/oUvo/<|Va|btwHw3+azT-K3@aNaGObqyw*yzwzw9zX+1=IqzbbbPKZv/bDumpCOKzjU>aL2pxjb2CF0Qaq0Yazb6bZa+1<3N;qE/u1bEa+b/>YJfv<HLv6b\\\"\\\",2):f(\\\"\\\"{b>ugfvxoPQaNz-/X:Dahy6u+R?\\\"\\\",2):f(\\\"\\\"}+o=*w\\\"\\\",2):f(\\\"\\\"}=p,bl*Y67bvozbkk2+.6c(dzbVaPacc+hdDt?>,bqeb>aub6+37LxY/L/hb5.,bhyz|5Aqr\\\"\\\",2):f(\\\"\\\"{p1A=\\\"\\\",2):f(\\\"\\\"{X53bayH/:Celmbyb<7ru.bmbgSBBjUEvF<v36<iQcbMG-b16?a156b\\\"\\\",2):f(\\\"\\\"}bWadGJWNaaI.G@aEE.b2phb=49:XajbZ=H\\\"\\\",2):f(\\\"\\\"{Y<=12u+bhrlb7b37FajbWaAsibyxzqn\\\"\\\",2):f(\\\"\\\"}|O*bTxebluyu5vRTG.Z3ab-=cbo\\\"\\\",2):f(\\\"\\\"}juH|O0C3\\\"\\\",2):f(\\\"\\\"}b|b"));
$write("%s",("JF\\\"\\\",2):f(\\\"\\\"}bZVV;lbWDxVuq31+h>DY3Dapp=xaXAaI762mA*YYa@Aj4U,.xMnK|9wV+=EZP,bXPX<y;SPTaZXko.6csdDzfo-o1|VZEPdD.Sl\\\"\\\",2):f(\\\"\\\"}+S:U.B/C>SKoYqlbZ>>G-q.bV++oIqWCdu4tntbWjbbEk.6qEazI,bGyL-1Q.h>xnoY3Thz?p+EP-1Da=ENG?RThz?Da-EDa>GDa.F+eCyp6|6yb9TVn>GV+?tV+wbDa=q@Wjb|p9mMM6bS|@WRo;OUaJvHnmzSaUtM8b4-bVa,bs/:Bco2bTa3v:BcoY+Fa,baok+DNA\\\"\\\",2):f(\\\"\\\"}Roow9F0xV+.Fro*ZXa-bY3z1H:2rSaZAA\\\"\\\",2):f(\\\"\\\"}koYJVnTNV+tbQN/2/LS3Y37vzI9d7cEagoVng0.\\\"\\\",2):f(\\\"\\\"{rOV+c7.tbo1Albz;8Nq\\\"\\\",2):f(\\\"\\\"{-FpLufTaS3/L3b.q>aWq7bS|\\\"\\\",2):f(\\\"\\\"}w\\\"\\\",2):f(\\\"\\\"}N7bubWJRaVn.qjbWJ.bV+.qjbbrAaax2b7bubbr>ue23bF\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"{4.z@Wjb@a5bNakb1EFaTa>+?acrCsOC=hMpF*\\\"\\\",2):f(\\\"\\\"}U\\\"\\\",2):f(\\\"\\\"}rDalX8L7bV-fD?eb+mLDapBTx/pRaDMBM2z@MPzDaNg<M:UN-aM:U?atXO7=4PaDamb9N>4cObbhb-ko3au"));
$write("%s",("aDatXWpzM\\\"\\\",2):f(\\\"\\\"}UPk>xBJxz=p\\\"\\\",2):f(\\\"\\\"}3e#aJ=Lo0p0TDansduhb7*N-s=0pPkDaLn(6c;cCaY|VaFa/qeb?aDas*qwP0vHhug,R3ZaFaQowbMzjbh9|bSaDaxbxpFyzDEajbgVC\\\"\\\",2):f(\\\"\\\"}rqmtc\\\"\\\",2):f(\\\"\\\"{|bTvEZ,oe6tL;<PpB3AoACDaG.1K>=bACa7v+bCa9bhbZBguybCMjw=a@aDazz5rY*YFQtsqJF<pFrHoVav?/bOamy:-Oq+b<akb*oiL6+<a:CHp1pC|Vzvbebdml8BWOkJ9YBTahzfzhbot4p4v34zw6b+b(4a%a9xAS0bh-h-lrZBcbBG?aybo/OGV0Byi-#3aJdeb\\\"\\\",2):f(\\\"\\\"{oF1Cyj0F1CtXCq0jbL;Q7/l0RuV.Rl:.JyNA5lTxqitioF|K|L-u>ThRA4.pUNp=-ub>ajowo++-o4u3zL-+@XatYL-Da@aThzGZa7bctv*qGDalzPRurxMtbYan.hybU@a?>zb|-+d2*ub9>xb3?-iQastlX+hVaVaWOc@bbq*LWxbAqEaub;Lgbeb+b/yYanzbq2b7Dkb/V>\\\"\\\",2):f(\\\"\\\"}xbI+P8Z4Xa2=YIUg7E8\\\"\\\",2):f(\\\"\\\"{Th<xqsz|1;8b-bDKlbY/+XGyxbtXs=GLrp|YgB2vo8DaPrsj?zcb||=A.QBW\\\"\\\",2):f(\\\"\\\"{rmb\\\"\\\",2):f(\\\"\\\"{Z7stg;B9mn\\\"\\"));
$write("%s",("\",2):f(\\\"\\\"}Nr3C5r?DtbfoK,@BGw9pw7:C[9cxd<a-rzc,S*S,0YT67xbdbk=<GC0DH1|S3CqS3E3Pasj?z,biQj@Pyy<Fa\\\"\\\",2):f(\\\"\\\"{b8b.t?a-.;|QY?o|bwSPRTaZ*Nakb,*Pkdw3bhxgb*xmbm,a+NPXajHJ;3z,0m\\\"\\\",2):f(\\\"\\\"{L?E1LEThMP1|iL32DQi/OX<GCu.\\\"\\\",2):f(\\\"\\\"{xMkbMMYJn\\\"\\\",2):f(\\\"\\\"}yll6ojyz=a@vhb*vnHIqZa9bXaj\\\"\\\",2):f(\\\"\\\"}Lqs/7bib.1yU\\\"\\\",2):f(\\\"\\\"{YWN-b\\\"\\\",2):f(\\\"\\\"{oU4:u9pRL9wBoub<:q4Va7bcbwGcx8rJzgbistCqr>q/i+\\\"\\\",2):f(\\\"\\\"{tGK9,qux.22I1/l*\\\"\\\",2):f(\\\"\\\"{E+b<aebdLUaS3VU~6cnb0XZu/w26MpTaWyk=C|Zub1MsB2YfU\\\"\\\",2):f(\\\"\\\"}BzG\\\"\\\",2):f(\\\"\\\"}yb<ars6|@z<HOqV=<V<oupeb?aWTZqY=fM;|@a0,IvO7.4D-MPvb=qkx=q\\\"\\\",2):f(\\\"\\\"{*abY-Hh+3e;a<a?=0xBaGao>Gy:WO03A-*xvZ>,M3x|-QOOO.K++Raf@\\\"\\\",2):f(\\\"\\\"}u3Ia-G1yuw3albxbc2fuYfw7XyrhAaGa/G*2H2D-nyJ4z|8?I+RaC\\\"\\\",2):f(\\\"\\\"}AqiSDaw=z0ntlt2*FrK|4vE*g|a+f-atUaB"));
$write("%s",("VtbgrOaE+@\\\"\\\",2):f(\\\"\\\"}5yOa\\\"\\\",2):f(\\\"\\\"{Ys0.uPtn6cYaXadbev5L6Ru+Y6gB4vE*Oakk-b8V9J\\\"\\\",2):f(\\\"\\\"}Ac:dzjoQ*\\\"\\\",2):f(\\\"\\\"{w2bPa/|Sa/H.b=a>s3i*qi;jb\\\"\\\",2):f(\\\"\\\"{wYsPaFZRn?aQ*\\\"\\\",2):f(\\\"\\\"{wo/)3g\\\"\\\",2):f(\\\"\\\"}a8+ZnBzPNdb>aE+pze4fM0rl^127^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^32^[2fha\\\"\\\",2):f(\\\"\\\"})3(f\\\"\\\",2):f(\\\"\\\"{#v3rga(f;)0,73-Ubb1p+oO+fCJ94X3+1+Qa,d/H1bG1JK=a.rj@uv+0K*qg\\\"\\\",2):f(\\\"\\\"}b;5d>qpHP=>Ea8bJ<ht7A.y6bs/Wqn+9p9>S:uwxPVjcb3-mx37X+18u-379D/b80*b<a6bbY9.2b9p12Y3b2ybkB0T5Az|wkVag/X19mOn3bjsb><aPI+1ur7b/7cbdd4du,x*bwri/OXnF|<f2-b?a|bTh<x:vPIG4Aa.qZ/RZ>a-i7+5+gtXaAa7swz\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"{v8:NdtPabb?ag\\\"\\\",2):f(\\\"\\\"{A\\\"\\\",2):f(\\\"\\\"}-oUa9@pr.bbME1Vmc2.Lox3zK3yb-bVavbaY7ERoxpZAvbuwPa-bV0b>V"));
$write("%s",("mc2jb4byu;-tQVad<7A3DTa=1m,\\\"\\\",2):f(\\\"\\\"}b<rMn7Km0d1XQ41K6U6k7M|urhbuIP6K9yu:kl\\\"\\\",2):f(\\\"\\\"}G4ZaZs9N@aHLvs\\\"\\\",2):f(\\\"\\\"{b>aP=4+jyqOXC?aP6n>PaVa:h;|Vab3,;1pybL0e3TLy=aqa+dBoe44Q2?.Ob4U6:Rd;b31It2n+PEm7D6@aj7H|Vy?a.UJ+fzQaw6|b7b+8Aa,bpRhMnsZanqmbGR\\\"\\\",2):f(\\\"\\\"}CjR|6E.C8a*.K,qux\\\"\\\",2):f(\\\"\\\"}9VacbTambtCs-3bXwdbfbgy-d9qQaS2pYL73@5b5r=aERdt2\\\"\\\",2):f(\\\"\\\"{OEQnCa-bz\\\"\\\",2):f(\\\"\\\"{uxZaOEh4a5bJ*>:bWPJS+BaS3:x|mZ|6545U5wu.rQafDib*btb.@V4GzxW8Rzs7AU5W*PRF0fbUxbLpR@Q.CeL@atlJzSa9@==9p7X9bK6EaQa?r?vNpLR1q:oSoInuyWTmb|-0rTxLoXT=F?DDdydabTNo\\\"\\\",2):f(\\\"\\\"}TN|-dbw4:oSok50<Dnc2gVg=Sabbxb<a9b6beb.1tG>\\\"\\\",2):f(\\\"\\\"}yWhWZqp?Zqp?6bLzMp@,\\\"\\\",2):f(\\\"\\\"{ys/*p2=ex=CNa?a:5W95GXi5bNatbQv\\\"\\\",2):f(\\\"\\\"{bjbWyS=\\\"\\\",2):f(\\\"\\\"{*<v<Q\\\"\\\",2):f(\\\"\\\"{Y@a4w;0-bi.\\\"\\\",2):f(\\\"\\\"{tlo"));
$write("%s",("3b><>>X+tjfb>ywssg><okthkb?3U6J<2oY4mFhyMfL?vs,xlo3bntNN2u3K9Nv-R6CuVanQFpGzntkb7b.bhU@YRa\\\"\\\",2):f(\\\"\\\"{bL?g/Aamz3K9Nfr@abbp-=xH2.UX39N/bvb\\\"\\\",2):f(\\\"\\\"}xmFTL+v>a7px7GaPSab+\\\"\\\",2):f(\\\"\\\"}Dq41D4Rd~d||b0LO\\\"\\\",2):f(\\\"\\\"}bkZCnWaB-M6ZaybUO:-NaiH/t1E<t<ai\\\"\\\",2):f(\\\"\\\"{g.Nyy1n\\\"\\\",2):f(\\\"\\\"}EzRaXy,tFp>aJh74ybs*ybPzqpib9paVz*+b3Ief>P<>\\\"\\\",2):f(\\\"\\\"}b>a:MCtDPRa5=OXF,At.-0xBaa3VjpUiLU4<a=sybNatw,b.bPr\\\"\\\",2):f(\\\"\\\"{b;sSr-kjr\\\"\\\",2):f(\\\"\\\"{b@z@?\\\"\\\",2):f(\\\"\\\"{b|qIDvlu>Na*b@a5bFadoq0.7WMtJ,0-bx0gbcxPB-=f7+bVZ0C:go=j9Fv?|>+3t-t1=>\\\"\\\",2):f(\\\"\\\"}CXOaT7m\\\"\\\",2):f(\\\"\\\"{/>nH|<>tns@AOtFa9wgbdb2XTajR;sP8<*Va.KOa\\\"\\\",2):f(\\\"\\\"{b,FwLw;jr(6cpdib3+HqzwHw?a1bD+41s1;r.b-b;|:xiBNpysRagB..urDU2+Zqys8wR6FYwLRahb,Nq6AqctL/wb>5l6GvWqwxu\\\"\\\",2):f(\\\"\\\"}M4wk@AOt;|ub,AQaDaiFzbgOzbzb"));
$write("%s",("nZ9vwLdbfb97FIDI=pR-Z9dypsQ2NGZ<GM\\\"\\\",2):f(\\\"\\\"}b022?KnBBH2cbGzQvpHGGdz5rL?=A\\\"\\\",2):f(\\\"\\\"{b4v2Q=xdbAJ4zebN=VaAJ6D;se4e08q<a04SP.zmb5b.zrxebjwWvR6:DhU-Vtzc@ebBsnHq,=CY*ebdLER52Onp@4Q2Q=x|RicaZmx4a^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'c0,/b\\\"\\\",2):f(\\\"\\\"{b-E>N.t<>\\\"\\\",2):f(\\\"\\\"{rs-?t:y1bd|8MYRotmtktZa7bhb.x2bYvp\\\"\\\",2):f(\\\"\\\"{f8eqKW-dhU=V1tebjbxbVUbb48OnZ|Kvtfbb>Nq*6b+b@Jyb\\\"\\\",2):f(\\\"\\\"{bjbis.v3K.bwvybx=z\\\"\\\",2):f(\\\"\\\"{*vHqr:JxX:jyGAlb6\\\"\\\",2):f(\\\"\\\"}EzyOysLEnHw;+F6gbb6b\\\"\\\",2):f(\\\"\\\"{bCaKH-dGR32mz;su:9yB+gbOacJfhGamVc=6b<Kyv9w7wZkWPhbOH(ba7kIvZIvba7ZI.da,43?4[ha(f;)59"));
$write("%s",("4A4.ia(ntnirpnt41da652t4.ba)T5[97[97[v3lqa:4*4>Qgb;O@va->og3a3aRopUcrOXF,c0Eau6GAKG.,jb3bTxM;QYW@\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"{Y<?aIuc>n8>Ac;aJo*b?acz-ijr\\\"\\\",2):f(\\\"\\\"}rSa:vq\\\"\\\",2):f(\\\"\\\"{c7I<QaQx/9@a|brrLF3ka\\\"\\\",2):f(\\\"\\\"}eW4Rvb.L\\\"\\\",2):f(\\\"\\\"}bh>i3c9cC03?hQbW5b=aD*euvg*5Cao/tMkkS/zbQx7tquou*.WaTBNWSa>FnyJxY4CaCaSaTO2z4z+bmb||.r\\\"\\\",2):f(\\\"\\\"{3fLvb2sZa@a5tw23oOaKo62S.rxvudycbvHNawxeb>aYvU+\\\"\\\",2):f(\\\"\\\"{31@abM>F;@s>qxbvb8bZak=luA7/.=7>7lro\\\"\\\",2):f(\\\"\\\"}0rjH,vTxArvb6.mIYCYT67lS>17xV4?aFJ>,L76eqg=;HIAaWah.w7vbVa><Ks&6cdbYayb\\\"\\\",2):f(\\\"\\\"{bXnfojbcrlXS6XahG9pr@GLNy-F?3L?7bb7vl|bqgH|HdH/hDiX1@i/7bib\\\"\\\",2):f(\\\"\\\"}bTBgyboFH-bZq;81Y>a>z6bWvg5aic7v@:q>pou:K9+y\\\"\\\",2):f(\\\"\\\"}b3bIv=aF*7br6zbj3em\\\"\\\",2):f(\\\"\\\"{*ffh/<z>P12Y3\\\"\\\",2):f(\\\"\\\"}bp@LEWT98hb?W/b@QS\\\"\\"));
$write("%s",("\",2):f(\\\"\\\"{>G?XO=YJ8bCi::ffw5kb1zGyubIBS=K6In\\\"\\\",2):f(\\\"\\\"{DGL.uarXs7*=qkxs/ub3i\\\"\\\",2):f(\\\"\\\"{uCn0CiQpUxVA\\\"\\\",2):f(\\\"\\\"}V,bD,Yb1JT<r80h/fbs1;|Jn1bdyOXnFWz+\\\"\\\",2):f(\\\"\\\"{OaOGvb?;x6c$akkm;8Pw-9pn+Ta/b=aD6;EZ>r;p;Ta/$Y[$YbYc=aVaQaxy-84b5\\\"\\\",2):f(\\\"\\\"}pz+ed/6.H8GLQ2G8cbjbqgD;@t.b?==\\\"\\\",2):f(\\\"\\\"{G>b.jtbb,b1DxqY62TWa9P:D@s2Ubbjb70Vm|+k|Uab.S|Rtib\\\"\\\",2):f(\\\"\\\"}<5bWaZhQ*qgD;TaQ6SaWa3b964;=a|+f.lKcG@a\\\"\\\",2):f(\\\"\\\"{X/QzrJ5NEtbfcVa1;/bRaoKjbxbzbzbRaTa8bcdE\\\"\\\",2):f(\\\"\\\"}Salbxb/QBwxM18Wz?P70ab|:Y/PaJ+j76bC\\\"\\\",2):f(\\\"\\\"}y9Eu0p9rJ+tCu.l3M<:g.ExIAqabq5FLRAc7c4d/fu?L<IitdFcZa.u.|Q-O-/p|bCuDadD0b*pbvupc27rc7NaL=UaxVfhRa1bx=LRTzsYOa?=\\\"\\\",2):f(\\\"\\\"{7XyVne>PkMyYarsi>L7Vast3B0,:q?=sm97hbj9Yayg\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"{o9ry6PT-6P/b3Xc7,dq6M><:A4R>Z\\\"\\\",2):f(\\\"\\"));
$write("%s",("\"}KF?Dr1x3\\\"\\\",2):f(\\\"\\\"}bZ<|<P==aq|>P<af.A?mA1u+0b?S+c2.vkQQn:sDaHC9bhb3+hc|m,bbb<G,bkrVa18,/PKZ3Z>Z3nh5tLWWaX*m7=amDy0C8T6sowqx75yjvPa5vZPlCjbSr-kIuVaV/kbWz9AeNb+b>DNZbV\\\"\\\",2):f(\\\"\\\"}I6b/EzvGrg,>aWaw7+biLUa@aOae9;t-bpUJFlbot<|T@Wac:OawP=SF\\\"\\\",2):f(\\\"\\\"{Ua;=ikVa9bpU=a>5AtPKybQrR6-2@u<:mA2bBW.b=akb+yF;kql*e4Vagb@uVaJ=L=9bz\\\"\\\",2):f(\\\"\\\"{E>31;0,o9kfFmA|=Wz\\\"\\\",2):f(\\\"\\\"{rzAeb4OaqaebbLUL3bwL*bCagbc5avbPkZ9g.5y+8sFYso9fr:-LR9pRyLt/bkYa*08EaFt/@C8q@ibcrlX|-Z3j@f/As,bmb*3ZBgudbbboDgbY/y9Dar,:vAAhuWadbTr.>ibe|<>9Ze$d7-/t-tO@E.eyJ5hbVz;0mt-/j6E2-vebW<cbTrRv.64QZWH29bCuQa+b:D8->aF,AtFnlt?>Aw=pcx?aD6jb?aIufhp@MU=1BwmNqw<T9N1bvbhq?3YSF*ntltRaZaTsUam0yuHD9o\\\"\\\",2):f(\\\"\\\"{LKEaAm.TrKocwBy6bCu7b5b4+?98bzw:vAAdLUaAq\\\"\\\",2):f(\\\"\\\"{JYnm,\\\"\\\",2):f(\\\"\\\"}bJ0P0cbEaRvFTx-yl3"));
$write("%s",("+cbEa5@Vfm.cbGzm\\\"\\\",2):f(\\\"\\\"{*I54GaPShqL<4QmF@v->Kv-bhb?aiy*bAA2XmbdbcbA:m\\\"\\\",2):f(\\\"\\\"{ibw=GCgocbD?Jo+bYaF|05U.,6c|dWnThlP6g|v\\\"\\\",2):f(\\\"\\\"{=BBmbub?|yOxbyU7sAaFyRayb<aebjb\\\"\\\",2):f(\\\"\\\"{E8b+8+b:pM?z8Za,v-yMq4RCaA/xb9>R\\\"\\\",2):f(\\\"\\\"{Thnyb-=axb*31y?/\\\"\\\",2):f(\\\"\\\"{bxD2D1E.vK\\\"\\\",2):f(\\\"\\\"{9>Wa1@4Q+b<E,EEaQYTh/YiFcw4wJ+tj.00bgYcbK<y+Nt;ECtUtwz>afFz+>rSzUiF\\\"\\\",2):f(\\\"\\\"{QaY4>a?o7HMzWaxsVg*bwbWClbVm>avLL;HJOGhQ:MLvxR7sRvLvBa<EHCw;Yy,tH7rqvlPHy=iFbbXaJ=GOLv5+fE7b>:-/v;=1BwU5*bRamNqwCaDD&6c,d.4WBy=osybF\\\"\\\",2):f(\\\"\\\"{FacbjbfT0rCiaxkbZ*.2bb-Say*32ohVbdf.EaxbBzPNAaxVSB-k1Eb7S3<a?=rON=VaFalovbhbkoUavgU17f8EG1\\\"\\\",2):f(\\\"\\\"{;hbRvGK?=ebBa<4bABaV\\\"\\\",2):f(\\\"\\\"}GKu.GzCa.diG.dytbANA@VfwhblA?aM<7b.bLp5G1bSa=a/tfbRacb.bwzlbubxH:vSabAxw?aEa@asE,LBaAa<4zdUafbBa+9JVub"));
$write("%s",("SaCH.b@\\\"\\\",2):f(\\\"\\\"}k.31+zE,hrfbBaQwXqGKu.oubb5GBwiMXq\\\"\\\",2):f(\\\"\\\"{bB4Sch\\\"\\\",2):f(\\\"\\\"{AUB4bAxwN@.r+\\\"\\\",2):f(\\\"\\\"{<4>.zA2X\\\"\\\",2):f(\\\"\\\"{>06aEaQa>;y/-/ubxHV49pCaV49p=yU6,p\\\"\\\",2):f(\\\"\\\"{srq9bw-r1E8Ta5b?HTajRLpjRLpThat,23by3aQaE8F0m,cbs*l@Lv0bkO:x+bbbibAwEaSPldOaRwv?yb=\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"{rvx1\\\"\\\",2):f(\\\"\\\"{JYNatbxVjub7AGG0@rx=1s94I7c7c:b;hwvdb@At2KsASS2INc=g/@,g/N1g/Rn;y|:>.gB2XTaTh?l;sfhJ8jwyuPa-bAG7J+h31+8FacbtC1sf/kFibub*.eczY,0z3dT7f5\\\"\\\",2):f(\\\"\\\"}ApYSC|.xHpvb,NY/hb3b5bYa=CVaQ5,/rG70zLdqubXavlfbgb4Yo\\\"\\\",2):f(\\\"\\\"}nF=aQ/mb/b?vPqfbmr4i::Fptr/HN*-BMfaO7bhb.x\\\"\\\",2):f(\\\"\\\"}bv8y9r-+Fe0..E11s,bq\\\"\\\",2):f(\\\"\\\"{:vq\\\"\\\",2):f(\\\"\\\"{Mv+N>Nc2gVg=Sabbxb<a9b6bWvkbRqs=.KMMG1,;2,nqBOyv2InHG1,T5b:mwbTa0qQYU.mbo7+EQaPa;s0o28Q*V,/>vbDaCaK\\\"\\\",2):f(\\\"\\\"{"));
$write("%s",("eI\\\"\\\",2):f(\\\"\\\"{bX*oB3zFav9HUx-@?.x;4QazA>-a6to\\\"\\\",2):f(\\\"\\\"{Z\\\"\\\",2):f(\\\"\\\"{=vutbqx,3z;tL.oKHtG8b1?huHsh\\\"\\\",2):f(\\\"\\\"{QD?a>OEaGalIkTKvLO?\\\"\\\",2):f(\\\"\\\"}NxGxf\\\"\\\",2):f(\\\"\\\"{0,fb?LsR.OPE4i*@q<xBdXUx0bT1Txm2p2VqPafb?/\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"{Iuqv>4bb@\\\"\\\",2):f(\\\"\\\"}6bg.>a7t@\\\"\\\",2):f(\\\"\\\"}ZDRa:q7b=ay/RF.bZa=\\\"\\\",2):f(\\\"\\\"{D\\\"\\\",2):f(\\\"\\\"}xb,NyWUD2bmb;5,bhxVaAz7TW*R3Ca9,wbwb6bemj;>V4z0Oub<a,3C\\\"\\\",2):f(\\\"\\\"{X|q6H\\\"\\\",2):f(\\\"\\\"{j-Q6FJHw=5wbR3L<yw<atblbF0X<5qtb@aMrfuTa=aF+Kv9b<aJT0wgHvCW+wb0TFK-zdFe0m6MyNpHqtjwz|d;OfLF2EaAoGT4j5bkb5b.b-dVfAs|Uq6wb1bT-6p5=xbY-w5FUp\\\"\\\",2):f(\\\"\\\"{H:Ep=a\\\"\\\",2):f(\\\"\\\"{b,Ni*jQZHubmKwbZPAq?\\\"\\\",2):f(\\\"\\\"}G5\\\"\\\",2):f(\\\"\\\"}@-J\\\"\\\",2):f(\\\"\\\"{@sVRJF8+b\\\"\\\",2):f(\\\"\\\"{b2s?uO86.ubRyhbxI2bGu3oeciVGy-zWawx6Wo;3WEagy0Wcb.WEaPa402\\\"\\\""));
$write("%s",(",2):f(\\\"\\\"}vzLmzb9y,|\\\"\\\",2):f(\\\"\\\"}W\\\"\\\",2):f(\\\"\\\"{Wgb9khUFUE3mA+E9b.-:yewHs@07bN\\\\\\\"\\\"),\\\\n(\\\\\\\"\\\"34\\\"\\\",2):f(\\\"\\\"}YaB*=+7RWaMrjzgy8/Au>v1.iW*qkkZV3xzb+yPRjb<:QR3bxI.b90+=B:=@3:S,?><EKGq5YsRyzbAs=qpqVaV+kw0V;tUa/4G.b::DGG/b.zvbT,MM:Bwb2zh\\\"\\\",2):f(\\\"\\\"{7|zAR3BoMf|z5b;<u.WnI6Qvl3XU.*+<t.-bN.o:+Pm1tTKIf/Ao@aO|x+hqt.8J+bvbTaAoPkS3iqGae-:Dr.twld,bqOv*Q7\\\"\\\",2):f(\\\"\\\"}rLKSar35G0v7|tb0:CuAoEaXa=S:B6bu.Sa.1ib|LyqzzWBjbubut.U,;Sap?.o*yf/\\\"\\\",2):f(\\\"\\\"{Ef3UawrS6-rsuhbtbcro\\\"\\\",2):f(\\\"\\\"{CahUWzRaluax8=kbiUTP0iYae5jrB\\\"\\\",2):f(\\\"\\\"}PaGarPMKpRAox=GakSERn.l\\\"\\\",2):f(\\\"\\\"}Ga/*/\\\"\\\",2):f(\\\"\\\"{vbWg<|zbI-YyitL</>-rR<kb-bYaI70b9b5/M8ybitvrd?9bUL\\\"\\\",2):f(\\\"\\\"}ba9YRvbERHrY=Qaxq37Ca1@Qa;|.80ssjj8@B8Je5V?Qa.4G553/RG5-RY<+0V4BBCanFB:\\\"\\\",2):f(\\\"\\\"{r4bO7K?6.GIkbD,GFB6cO\\\"\\\",2"));
$write("%s",("):f(\\\"\\\"{J1bwbTNUtiw8r:+V/-IO|>2G1?v4+?yz+nQ6vyOVswr0b@RayUK5bR*E?c:+be+I6YIz\\\"\\\",2):f(\\\"\\\"{aQ=AxDxECrk3089pg,9qybOavo*b+bTL5i7J\\\"\\\",2):f(\\\"\\\"{f2*cwY<yzANqsY6*b1b6,5.aorwThpwO0P8CrFa\\\"\\\",2):f(\\\"\\\"}4T\\\"\\\",2):f(\\\"\\\"}PN8=\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"{Q\\\"\\\",2):f(\\\"\\\"{ko5bQrX52oi|KvSK41ub8bXs<@>AS?X,+=OsGa5O*NXaP8YqdPZt:<ubL<9>Xt8wB*mbFj-b/bkoxbVqz\\\"\\\",2):f(\\\"\\\"{G5j1n:N.\\\"\\\",2):f(\\\"\\\"}PI8Xa5bdbXaTv:x+8@a8*gs0bHC.bHJ\\\"\\\",2):f(\\\"\\\"{0abSrQruNBNGasO4+zqJ80OT7Patb-3X>t*U.3bUtxv4bl\\\"\\\",2):f(\\\"\\\"}fbeq>N-iIvjb-g>JMofqnr*qAqt*Pawru-kqmDcbUxCa7bqO<uYaEa8vBN+hl*Ya1bhbkbT+2b>a|pQqM;?rXa\\\"\\\",2):f(\\\"\\\"{/Ta?vZam\\\"\\\",2):f(\\\"\\\"}*k|-ubJhPsb.OLc:Wzwbkrhul\\\"\\\",2):f(\\\"\\\"}8bDa9pX3zolCFyEazb9bZa/7y+lbqsThT<.bPN:ohbK39p1bdL1brp*5YytLNEPaOa7b>@su1;Sa^127^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):"));
$write("%s",("f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^32^[2fha\\\"\\\",2):f(\\\"\\\"})3(f\\\"\\\",2):f(\\\"\\\"{#v3rga(f;)0,73-c1FaR-WIW@prWaVa>ofbSavb05*bfo:,P-+C/l13|@m:xN4bebf@w<WaRa56uqoD4*;qGyC\\\"\\\",2):f(\\\"\\\"{FaPa9p,bzb|tlozbJ3-1+u\\\"\\\",2):f(\\\"\\\"}bNG.?3w-ERzybmbLmebfbc50|=+Xa+8Ft1sTao.SK<vSKNaNaU.vDQDkbhMszNafbXnm\\\"\\\",2):f(\\\"\\\"{Oa0,Xy/>D8=jD@KDt|C/ZaUaH/ebg/urTn;LcbSaaOeq>a.b/1\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"{yt*II9Na0b@rG.Aai>1pEaYs1\\\"\\\",2):f(\\\"\\\"}98dbjD0b1zdb1blb6b16>a6bCGHClb8*fjTaFaHJwbS3qs7v32SB@B>a9b.bJ9XyabAqA.nr@axb1sxb>aPaMpUaY\\\"\\\",2):f(\\\"\\\"}h9M=FqN*nky;fb+N8Jfb=a-bV|D.LuzB4H*Lelqs|baA8*oMcbZa5+ubYa9bB9\\\"\\\",2):f(\\\"\\\"}bfbebh/L9N=*kbJ+hqGk3fzwtVaybRa+b.Eayc7B4sHBM*b<:?HgvHqYv0bvz8wDwbbgb/=m+7.NgYazq=\\\"\\\",2):f(\\\"\\\"{Oa.8CaE3D?x7lr1bxMME*MxMPaS/VmR|pMbb<wu.MtHq=a*bR|"));
$write("%s",("\\\"\\\",2):f(\\\"\\\"{rLw/bm-rxp?8bGKS\\\"\\\",2):f(\\\"\\\"{zb\\\"\\\",2):f(\\\"\\\"}bmK4v*bs*kb3rRn9B<a;o7tR3JqC=t|wbcbVl*b>,|swz?aMn9bvHj3|9Va8b4*,ut*q3wbo.7btj0biLOoNaVCn/yb.pcJubvbHhz1M8MojbFa:6jb2H*J,b3br6ApdmPpxbybj+wbY*-b9bPaEngCCaWp|EF+,bAs?CQazb<aAJQa:g.8\\\"\\\",2):f(\\\"\\\"}>.8fq@r3qtF0b-:EaebkFJd*.4bB4VaY/z6Bai/Lpi/31Fp;xf\\\"\\\",2):f(\\\"\\\"}K7836-Ba.bfxb7MB2uvz?r367bypwbt4tbTan.mrL*dbPaF3D3B3SoQoyIjzNrNoLoJox4ju3b5\\\"\\\",2):f(\\\"\\\"}zbIhgb+omx/9Kx:oXs|3Pr3o\\\"\\\",2):f(\\\"\\\"{|g0vb5y7bM4Y/V3nvEa>p/b/74wF17sacCo4bOa8uvbV-YA<ajb1btb4bgbq@6bo+kb?aubdblu=uqx5bM;6zs3inG5yBbswB2H3q+b>aBoGw5qJ.oD4/tb2/Q,7-iqvbm7W*rwSaSpdz5t3tJ8t*6I/b\\\"\\\",2):f(\\\"\\\"}>ub=pkbk|KH<:h-9b*dU3ABgb7I>o0qg9lbf3c4Wa4b?abbfxT8.7-rM8db05d>Qae:TaU:y9Yv94o+x4ubBaWa94s/=awbm;b1ThnG=\\\"\\\",2):f(\\\"\\\"{QoAa1bubhb2bOautQp|w\\\"\\\",2)"));
$write("%s",(":f(\\\"\\\"{=A4T;/7Th-?E.2\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}b=a.,Cscufxgb0sSanAayk@*;h@QttgUq3e.,zbEa9|,tIqib/tNA3b0qebttg=abO+qp2*dbf/Av+bgu@o7|e4q*Lud83FO.1Fdb;xPans:8D\\\"\\\",2):f(\\\"\\\"{S\\\"\\\",2):f(\\\"\\\"{V+DaRa?r:mSaCaZagbVj;49b;vbH?aGa3*iqS/ZaXai/b1a3<a@a9p<a+bb3Qq4z\\\"\\\",2):f(\\\"\\\"}6><H/U*Qa.:H-S/e9J@;<Ea,;Ta-b3kBqjb+.Aa;.1bNaEa96\\\"\\\",2):f(\\\"\\\"{|lb-2FaEtTBU6Ca1uqplbBq28/>4bTh9*u.B@pBB*V35be?YE?ad|3gR/U>KD.bCqNaxbjbJ96bv:ikN//uRaibq?7xVa5b*bD?/b;8?yt?z\\\"\\\",2):f(\\\"\\\"{p7;v@smbZa:\\\"\\\",2):f(\\\"\\\"{,tYv8b=@z3<a>a>.>xlbRwG\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{bV0P=fr=AA9Thq;9Bgb+bNawb5bc/w\\\"\\\",2):f(\\\"\\\"{t\\\"\\\",2):f(\\\"\\\"{p<33,D@avblbRaQaybT,avq62/\\\"\\\",2):f(\\\"\\\"{pMtUwlb>7>7UaybqxFr@a\\\"\\\",2):f(\\\"\\\"}bRa4boD8bmD3bJ00|mbTCkbRCL<.o+87@\\\"\\\",2):f(\\\"\\\"{80by8-:Hpvps>B27b<ERa2bjb\\\"\\\",2):f(\\\"\\\"}b"));
$write("%s",("b>vbfbYaIBabJ4M<\\\"\\\",2):f(\\\"\\\"{Cyhj|1BECzbTalbz6zzdb|b1DHCYqU3ftvbMz7v1ySacb=aj+<rmDybhb\\\"\\\",2):f(\\\"\\\"}b\\\"\\\",2):f(\\\"\\\"{byb6bPa=aAw7sNaaoSag004.*kb@t;<b>4+m|<:k-DaVao5\\\"\\\",2):f(\\\"\\\"{bM61@kbb>*btquwBq>aEa*bXaTnEa?ayrPa|bebc??C31L<+76b3bEagbJznz\\\"\\\",2):f(\\\"\\\"}-UamyWalz@a3kWacbCmxbv8xCy=*l*DbpuBz1wrurTa05RaE2PaSzJwtto\\\"\\\",2):f(\\\"\\\"}o57tDarxlbgcV+RaxbQa7:*br:>ab79bZhu-FaR3>a8bdyFpPvxbDsBs@sqgyh\\\"\\\",2):f(\\\"\\\"{b?>/Clb\\\"\\\",2):f(\\\"\\\"}b<ar6LfY*7*-bsuc:3bEB5bp?ypNaU5?=W\\\"\\\",2):f(\\\"\\\"{kooBxC7|Aa=aRaBa3bI+7bZtnjtbd?io1Bjb\\\"\\\",2):f(\\\"\\\"{bC|VaZ=1bWabo+b9py1,b=ptbAaqucuu.=aibF0Y3VaPwxo\\\"\\\",2):f(\\\"\\\"{b<a;3=aBa<alb\\\"\\\",2):f(\\\"\\\"{b,wBqdbz1/o2bO:N5XvG/Na|3/>ow@7yb.bdbYaizI?/bEaflAa<aA:@4/>x49qy=gBd0koc\\\"\\\",2):f(\\\"\\\"{wbPag|uhd0,bLxinN.c8Tuz@2lx@Oq@r9mU.<amb\\\"\\\",2):f(\\\"\\\"{;P->"));
$write("%s",("tzbOq2b8wFaw7-bp?O0n-WzQa6b@a90Razd?,h87bD*ZaCucbj*4<=AJ4gbld2s:|q4G.Mymodb7b5/Gae@|<upuh::7/mbx4CaGa/6Yvfb<aB4EwTzIqIxm|kkkq/>QaRvwx2w6>@?kv9h6|c\\\"\\\",2):f(\\\"\\\"{@<e*X81b-5<wUaf5k?:?,>e;1bs/+b0bdwT6/bNa7tb/2bd4g3.tdy7bzbI.Tqk,i,;v8bl\\\"\\\",2):f(\\\"\\\"}ts<qebw50bGiG1bb@40bzb8bM*cbsj\\\"\\\",2):f(\\\"\\\"}84\\\"\\\",2):f(\\\"\\\"}/ba;Aa>jzb\\\"\\\",2):f(\\\"\\\"}>7b7bv/p-M<N.o1F5O\\\"\\\",2):f(\\\"\\\"}l1/lz>R<Taj*rzx4G-Na\\\"\\\",2):f(\\\"\\\"{bS6f\\\"\\\",2):f(\\\"\\\"}N3Nad/gbi6g6-dThgx.6ub\\\"\\\",2):f(\\\"\\\"}oT-X27|C8\\\"\\\",2):f(\\\"\\\"}b,bx7ThIrmpI63>7yTh|8UaU*X5>amyDa6bEaBa\\\"\\\",2):f(\\\"\\\"{+=pRa5bd4E.<adbtsi?/tBa@28t@2d|wb\\\"\\\",2):f(\\\"\\\"{b?aXa=aJrab,tguZ4ewqu<\\\"\\\",2):f(\\\"\\\"}jb=+vs*0bbaz0b\\\"\\\",2):f(\\\"\\\"}wXv6z2b4zXig5k6px*xJ8C=hbj=abSaftAsUaAaBqibO34wXaC3J.+<huj|cjgy-bn47|vow;Tqeb?z1b/0Yakr=aB6ibq>wr<aqvzd>a4p/bwb9p<3"));
$write("%s",("Fp=h\\\"\\\",2):f(\\\"\\\"{oazXa::abQ;:.T-Taf*G5x>k1n<ZadbBaOaNa>y7bThI2@aBy/b*qb>6bjbqtGu32DaXy-b\\\"\\\",2):f(\\\"\\\"}rOa\\\"\\\",2):f(\\\"\\\"}bfh>tx=E1EpQaCt?=/bPkPa+bVaDalb,5?=0\\\"\\\",2):f(\\\"\\\"{D-3<u*8bGzIvfhNajb9bL7.blu>t@ay49mkbcxs07bSaB1woev.bZ4fb5vis\\\"\\\",2):f(\\\"\\\"{bYajy@a-bOaj=4e6bdbx<5bh=\\\"\\\",2):f(\\\"\\\"{bs11w>xfb5blb1.3b/\\\"\\\",2):f(\\\"\\\"{N7;sbbW|Yf,blbSa\\\"\\\",2):f(\\\"\\\"}bZ4<\\\"\\\",2):f(\\\"\\\"}.bG<9btuub\\\"\\\",2):f(\\\"\\\"{+tbcb/babBa|bojzwQa9rmbM3m0@8a9Pwabh\\\"\\\",2):f(\\\"\\\"}Ztib=a>jybvr<t@y9pM|/yY*O+SaH/S\\\"\\\",2):f(\\\"\\\"{Qxfb1;<a?aR-P-N-9pYwr3>.Twy9w\\\"\\\",2):f(\\\"\\\"{Exb8|,k:Wa\\\"\\\",2):f(\\\"\\\"{5n\\\"\\\",2):f(\\\"\\\"{u.6y<aXa>+,d@rSxw/y0w03ky1|fdbV7T7bb7wBarwxbYaUa3bzrtbG0SwNoxbl,/y\\\"\\\",2):f(\\\"\\\"}+\\\"\\\",2):f(\\\"\\\"{3z./y@a+b97/h.x1;Bs>0qwrxF\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"{7C88bEan+?a=\\\"\\\",2):f(\\\"\\\"{m;\\\"\\"));
$write("%s",("\",2):f(\\\"\\\"{bf2=akw>.vb>a9p|1TaSaVas2,qqw8bq/>ab;8b:x-5xbbb+yBtqu5b5\\\"\\\",2):f(\\\"\\\"}i8s0J1k/8tBaTa6b7|c:8b9bV-X1VaL:96=\\\"\\\",2):f(\\\"\\\"{Dw+beb3b:vq4kkjt4bEa0bAa\\\"\\\",2):f(\\\"\\\"}|eb0wBaz|4b5bQacb<rz19b2btgywXawrr3lbNrTatbJhcbqpK4lb8oc\\\"\\\",2):f(\\\"\\\"{?87bccw\\\"\\\",2):f(\\\"\\\"}EaSww\\\"\\\",2):f(\\\"\\\"{Q.03w\\\"\\\",2):f(\\\"\\\"{D5Z7OavuZ4BoYuW\\\"\\\",2):f(\\\"\\\"{-bAa|bGaN|k9V*3bq9yr+3jv/yXaUa1bF8RambTa9p\\\"\\\",2):f(\\\"\\\"{b2bRvokabA*FaCaVarqEas1i0+1z3<u.7J8=\\\"\\\",2):f(\\\"\\\"{m|>0\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"}i5\\\"\\\",2):f(\\\"\\\"{b2tqp*bN/suJtlbq+vb7bru,vwbR\\\"\\\",2):f(\\\"\\\"{jdlbP\\\"\\\",2):f(\\\"\\\"{Ranq*wt*E*vb;-C*n..bjb-09bS|4tTaj,bbZt=a,/Awc*Ca|wz/LwP89pR-ybgbj0EaP-mpkbyb4bybdb.bOaWa2b?3TauoG3quYaXaSp/b-0Mv4b-p+bwbWaWaFa2*VaxbJ1\\\"\\\",2):f(\\\"\\\"}bJd9pWa9bO+++\\\"\\\",2):f(\\\"\\\"{sSatbQtib6bxw|bYs/4Cu.1=aS*=^12"));
$write("%s",("7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^32^[2fha\\\"\\\",2):f(\\\"\\\"})3(f\\\"\\\",2):f(\\\"\\\"{#v3rga(f;)0,73-c1a3b.\\\"\\\",2):f(\\\"\\\"{Dr<|inw\\\"\\\",2):f(\\\"\\\"{AxE5CxB5luBaj\\\"\\\",2):f(\\\"\\\"{YaBa4b9zth.b1vNa5bB/kbkbV0db,tV/hbq6A79bEpyb\\\"\\\",2):f(\\\"\\\"}b8bkbAq8bIvlwgb,tn\\\"\\\",2):f(\\\"\\\"}Dwqwg02bSwDcgfOa9pj\\\"\\\",2):f(\\\"\\\"{*bSauoiq8t@a\\\"\\\",2):f(\\\"\\\"}+nh/bVaEa66mdVqF6B6Xamb@aSarxM,WaSaZ3?a7bM,@t2bkb>,H*|b@5ro6|RaAaFa/bSaQaEaAaVa0rvbGa;/4bhrLm6yEaS\\\"\\\",2):f(\\\"\\\"{Tab.c4/p96y0f.psVaTa>\\\"\\\",2):f(\\\"\\\"{Z3@ambGgQaNaXaTht-wbPw+oEu+bWa0bb+Sa<|ab@a5\\\"\\\",2):f(\\\"\\\"}kbkk*yjbTaltqx7-tb\\\"\\\",2):f(\\\"\\\"}bCa=ahbBakq..\\\"\\\",2):f(\\\"\\\"}bUao55i9bcbgbwbd4>+AaTaU4Ba0byu3z3ompfb,v*bw\\\"\\\",2):f(\\\"\\\"{C523Uu/3u\\\"\\\",2):f(\\\"\\\"{x\\\"\\\",2):f(\\\"\\\"{43RaVaGiPa0b1|QaC0Rv<hcz7bbbutf"));
$write("%s",("b1q\\\"\\\",2):f(\\\"\\\"{bmb=+Y|fbtb@/ybpqqxzb4tn+*yeb|y7tS/VaYaVa.r@a*w1bn+lbmpy\\\"\\\",2):f(\\\"\\\"}H|+s\\\"\\\",2):f(\\\"\\\"}bYa+-dbgu,b=amb4ju3ab*bOn3xZt6p|rV2gb0w:wjrAaW2tthbwbHvi/BscbkbAaz2hb@acb4bTayb<vtbEt9pz0?a1wcdNaybZaPrf.\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"{0bNp.1hb-b6+PaYaa*YuXacjj||blz9\\\"\\\",2):f(\\\"\\\"}Tqs0Oo:gabm.DaSapx\\\"\\\",2):f(\\\"\\\"{bubUaEa\\\"\\\",2):f(\\\"\\\"{tSa>a7b*d8bxbKnwbhb=qf\\\"\\\",2):f(\\\"\\\"}Xa*bnz9|Wa?aduN*fbab8b,q4bDaXnc1@a0bltabybm|iqDa>yN.K\\\"\\\",2):f(\\\"\\\"}i1gnz,M.n1LuVoabwbMteb8/@a/b5bibib4jmbluYu4bXa,/s*MqgbTrlb,b8b+d7-7b0bRa;|PkFa8b:2jrUgAz8b=pK+Babu+bZtohTazb4bRaMs/bZax|ybvb7-Vqhbp+Qay+zb>a02zdybz-@ad|jb+bu*0b<a*bFa4bWagbZat.rs<aZqE1Daf2/byb1bprmbM,E\\\"\\\",2):f(\\\"\\\"{nzYaKp,wQampc0a0stDvQrgbCaC1gbfbhb*.5bubB1wqdb4b+.H0g15b1oNa<aEpR|abst@-1bOa,b2b>r.yZnEsV/vbRa.bwb*b"));
$write("%s",("/b>a:-vbkbcblbr1U.\\\"\\\",2):f(\\\"\\\"}+Fa3blbcr8bYyevhbF0lbfb2w|b<wQalbtb0bdjw\\\"\\\",2):f(\\\"\\\"{*,P\\\"\\\",2):f(\\\"\\\"}/lM\\\"\\\",2):f(\\\"\\\"}N.\\\"\\\",2):f(\\\"\\\"{,P.WzSam0Bak07bab4\\\"\\\",2):f(\\\"\\\"}kkX+*pK0YaD*QpNvD0>jdb?a6+lbOqh,|b*.hb,bFag0.bububq04\\\"\\\",2):f(\\\"\\\"}Saxbd0b0eb4\\\"\\\",2):f(\\\"\\\"}Caxb|bH||p5b8r+oRafb>aWzTa4b6b0b>jlzxbVaAafbkrJh4plrPa\\\"\\\",2):f(\\\"\\\"{dtbS/.ofu5bPt.bebxbNv6blb0b|b=a=a4r8b2b4p.v9p\\\"\\\",2):f(\\\"\\\"{dzwiblufbJr<\\\"\\\",2):f(\\\"\\\"{sj1.*bmb<pYuAaabv|UzRa3b,bcbFnAa@s\\\"\\\",2):f(\\\"\\\"{|ThLsLo|++babDaubWafjbb1bj-k|F|lbWaZt\\\"\\\",2):f(\\\"\\\"}b8uPs6bXaTaIn@-Va/tZalbAan+vbOa9b3zX\\\"\\\",2):f(\\\"\\\"{LqbqlbUa4bYaSa\\\"\\\",2):f(\\\"\\\"{bVm@ar\\\"\\\",2):f(\\\"\\\"}G-xvAsjz2s7bikfbLuR\\\"\\\",2):f(\\\"\\\"}L.IbJ\\\"\\\",2):f(\\\"\\\"}hp\\\"\\\",2):f(\\\"\\\"},Da3b/b>\\\"\\\",2):f(\\\"\\\"}jbu.3bWaos-r0br,Hpwbp\\\"\\\",2):f(\\\"\\\"{DqvbUaz.l"));
$write("%s",("+ay,byb?a@s\\\"\\\",2):f(\\\"\\\"{wPa=\\\"\\\",2):f(\\\"\\\"{/b.bbbmdgb\\\"\\\",2):f(\\\"\\\"}bGz?z=zPa;tB*n.crzbNas*@rTz9xbbmbcbAa@aWa=aSa.bRacuE\\\"\\\",2):f(\\\"\\\"}0-3bTh\\\"\\\",2):f(\\\"\\\"{-Va4bOk1b1bkb.|Oadb\\\"\\\",2):f(\\\"\\\"{bOahbPazbW,+bXaWamb6bbcThHtTaCa2bScRa<apubq=a@,ub\\\"\\\",2):f(\\\"\\\"}bwb?a3gibCa0r@aabcbj\\\"\\\",2):f(\\\"\\\"}S,RaRa/b9pNaOaAaPaSaH\\\"\\\",2):f(\\\"\\\"{9p3b*bebqtdbx\\\"\\\",2):f(\\\"\\\"}|bNado|bdb\\\"\\\",2):f(\\\"\\\"{o1bUxTh-\\\"\\\",2):f(\\\"\\\"{<aAs.bib9kzbOa@,4bNaubcbH+fbRtmoZsVayq*b0b6,+bkbQa9b@aEaV\\\"\\\",2):f(\\\"\\\"}3tfb|bhbcdtb=aFabbHnO+2b,x@sUaCa?ambCwfb.b7tLu0ly,L\\\"\\\",2):f(\\\"\\\"}WuQ\\\"\\\",2):f(\\\"\\\"}I\\\"\\\",2):f(\\\"\\\"}gbYwbqjqXaybzbmbflJd.bfbOa0v9bhu2bDa\\\"\\\",2):f(\\\"\\\"{b*b9|2bzh0r6bUagbD\\\"\\\",2):f(\\\"\\\"}EaNa|b@ayh;\\\"\\\",2):f(\\\"\\\"{0bdbkwnuEnVambzbQtfq*b-b2bKwfbDa\\\"\\\",2):f(\\\"\\\"{+wxmbBaLxxuwbIzlb=q+bhbjbdbvbshAq"));
$write("%s",("Qp>aIufjQa5xRa8bOaBa9psjcrUa2bduuvn\\\"\\\",2):f(\\\"\\\"{Za/blbgbPaNambPaV|6t1yRaUaabdb\\\"\\\",2):f(\\\"\\\"}bgb.bWa7bkbGwwb/odbgyjb=\\\"\\\",2):f(\\\"\\\"{:wOagbDa5bhbibgb4vYa<a\\\"\\\",2):f(\\\"\\\"{bab4b7bWa:rysDaq*2vMr0blb-bt*PkTh|*db<aThlx*b=qzbZa?a9p*b*bOqTxXy2vjbOa3bdbUaPaNgCa;|\\\"\\\",2):f(\\\"\\\"{bUaZa0b0b5b\\\"\\\",2):f(\\\"\\\"}wUaXa<pab0obbbbUamw5xzbnwNzinjiN\\\"\\\",2):f(\\\"\\\"}fp2lhiRuw\\\"\\\",2):f(\\\"\\\"{PuVuv\\\"\\\",2):f(\\\"\\\"{jbeb<aQaBambkbSa3bkblbL|9p3xh\\\"\\\",2):f(\\\"\\\"{7h1pQ|jbgb0b7t\\\"\\\",2):f(\\\"\\\"}bvb5|;v7b4bQpabhsC|ay:ogu0bmb+b7b8bfrYvCa1zWaXa0bOaXa?vPaib\\\"\\\",2):f(\\\"\\\"{bib@awgibCtAu2babhb4bZa2b4bCaNa8bAaUaTh?wxbmbtbkb3bCa\\\"\\\",2):f(\\\"\\\"{r|bZnvb<aBoGq<v|bcbBaFa*bhycbAk.bVabb>aMsspPaFa?albLfibtv7hBaUambQa?a<aLnPapq-bwzWwXatg=\\\"\\\",2):f(\\\"\\\"{TaUa+b3bcbhcroEaJwXa7bCuKyYa>rYuxb\\\"\\\",2):f(\\\"\\\"}bbbD\\\"\\\",2"));
$write("%s",("):f(\\\"\\\"{abWa|bibPa\\\"\\\",2):f(\\\"\\\"{upxH\\\"\\\",2):f(\\\"\\\"{As*bTvEp3bPtVaOaPadb,b/bXv+s3bubZaub*pioubg\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"}b|z:yxbNa4b@aUa9p4bysAavbBa-bFawbin4aOus\\\"\\\",2):f(\\\"\\\"{QuBxDxdzbbzblbPaebTzBokbqxab,b<aPajw@ajbZaZngyKw>aebub?aCa*bYfCa9o6bDakwebSa4bpu1bab|bhoQovb-b>a\\\"\\\",2):f(\\\"\\\"{b9bxbtbLpts0bjbjsFa>pebtbmb9b\\\"\\\",2):f(\\\"\\\"}sVjfbibwbXaRakb6bcqlbebuv8b7b<y2bAaxw=a7t.dXa.bXaBySafb\\\"\\\",2):f(\\\"\\\"{rtbVa:wUa5bmb3bgykbOaRrfb3y1y/y4btg>a=aOajbCa|bhyLn*b>aabqvOtkb2bibcbibAadbAazbhbYaYtAa.bDaqhvu/bAambgbtb7bwx3bmbBvTa3bbqpu/b\\\"\\\",2):f(\\\"\\\"}sfb0bThTtRavu=a9pYaebIxayybAaXaabNwmb=aZaNngbWaexqt/x-x,bdbWabxLv5xAahbXaSaeb\\\"\\\",2):f(\\\"\\\"}bmbUa.bLuXr@xYrLu.lVrgs-b9p-b\\\"\\\",2):f(\\\"\\\"{b-babpt0b1uebAs8b,xqtNa1bPaNt>aZwYa=a4j7tAatbMtgb\\\"\\\",2):f(\\\"\\\"{bWa1bHqWaBabb.bkk9p"));
$write("%s",("+b6bdxex9p|b6b,bPsRaXaNaQaTaxbXawg=a4b8bmbYa0b*bOaqvlbibjbwblbXa4e*b=aYaRabb9pQa@s5bCaStwbRaabxbEaguQaFaOa*b7b\\\"\\\",2):f(\\\"\\\"{bicBavb/b9b=a5btbabtbbblqelYaFaCsxb9pwbZarsAtwbbbvb*bcr3rCaub5bZa1bjo/bkbebYadrab7bCrPakb/bGvvbZajbEakb+bUacb5bzb*b5rab0bXa\\\"\\\",2):f(\\\"\\\"}b/b-bZamb1b?agb6b/bWaYa,b*bTabbTrYaQatb\\\"\\\",2):f(\\\"\\\"{b/bcb6bmbfv5b/bbb4pSaJrIuYabbDa1qxs>pjreb7bfbEnBagbxbOa=agbubtb|bLuenSuNubngpZrLuesascsjndsucmbwbvu|buuXa2bBaybeb5bEa1b@a8bFq*bEaCaFtmb1t-becZawbJd?a*bItUaUaUtcb1b7bfj8bebXaDa1bBadbabvbSaubxb7bZa\\\\\\\"\\\"),\\\\n(\\\\\\\"\\\"=t8bbb0bcbbbYacbab/bttZaxb0bLpht9pBa8b/bBa@aub7btbdb*bAa9pSavskb9p9bvb,bRa7bNa.blbbbPahb1o3bYa/b\\\"\\\",2):f(\\\"\\\"}bOaCa0b?a3bTacbmbOacb1s.oebVa4jRa.qybfb8b0bubNa\\\"\\\",2):f(\\\"\\\"}bVatbfbwbibhbEaUajb8bFaibeb4b9pyblbTagbZbYqWa,b5qHrFr5bwbCa9pi"));
$write("%s",("bOa-suqWa>p|b5b,bWaCaebhb|bUazbro^127^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^32^[2fha\\\"\\\",2):f(\\\"\\\"})3(f\\\"\\\",2):f(\\\"\\\"{#v3rga(f;)0,73-,#kbzbtbysFa>azo4r2rfbUa8b.r,rjrhrVa.q9btbtbNa3b7bUa|bbbQaUaOaEaabzbWa=p3bebbbcb\\\"\\\",2):f(\\\"\\\"}bDainhidpWrepipcpinin<iWocbOa/bDakbFaioEa9pNgub9p\\\"\\\",2):f(\\\"\\\"}b6b7bdbwb2b0b@alb4bubabMo0bQoTa1bFa.bzoebgbQa1bBq8bUaQa.bNqQair?aabYaCaabLp|bTaYa-bsjFaSaPaco5bOaubQa\\\"\\\",2):f(\\\"\\\"{b.bUaSaYaubjbcb9bzbjbRazb2b.b1bVa6b?a6b>aOaib9b8b\\\"\\\",2):f(\\\"\\\"}b1bdb8b.b>ombWafbQa|b\\\"\\\",2):f(\\\"\\\"{qyq>aNa9p2b@aFa+bSaEaFa4gbq+oYa2b5bDaYawbvlgbNn\\\"\\\",2):f(\\\"\\\"{bPpmb4bjbNa<hkbRavbdbCambvbvb\\\"\\\",2):f(\\\"\\\"}bebmbibTadbrh9blb4gYaab|pjb4p?ecb/pFaDazbKpkbdb,ojb-bSawbjbhblbYaZa-bwpDaTa2b>p+dXabb\\\"\\\",2):f(\\\"\\\"}bxgGa"));
$write("%s",("FoPa4bvbcbwb=a,bZahb6bxbcb@atb>aRojb,b?akbibDaFa7b1bDawb7b\\\"\\\",2):f(\\\"\\\"}bylxo0bibvbjiYoZo*lXo*laphnjilnmnjikninNa\\\"\\\",2):f(\\\"\\\"}o6fjbPa,bukwbmbSaXaFa6bSahbThqbRa-bCaFa-b7bTaQaTnYacomb,bYa3o4o2o0o7b/bYagbib,bjbvbNahb/b1bebFajombXaZa\\\"\\\",2):f(\\\"\\\"{b=aTa\\\"\\\",2):f(\\\"\\\"{bwbEako1bUa>aFa|bWa\\\"\\\",2):f(\\\"\\\"{bdb-b4jeblbzb,bNa7bvbCaEahb<aCabb*bzhQaub*bWaQagbSa,bEa7b6bAaEaJl9nxn=mmmkmqnEfSmumsm/n;a@mtmrmSm?m<l\\\"\\\",2):f(\\\"\\\"}n-bJl6mCa;lPmwbicSm=ljmtnEaUl@mlm;lzmgmemin2l2lcn4afn9ahidn*lan-lji1l/b\\\"\\\",2):f(\\\"\\\"{f-a\\\"\\\",2):f(\\\"\\\"}hub/h8a7mDm\\\"\\\",2):f(\\\"\\\"{mIm:l9aEaOa@m>m/m8f:a-b@m=aAa-a0m*mCaUlYlym@a<a-b|e3m\\\"\\\",2):f(\\\"\\\"}mMlimXlOlMlKlpm|m:aCa|evm>aAajmTlOl9a8lPlAa?a>aFl|ehmulJlWlBa-aLlElCl*bvbtb/b-a+bId>lQl?lHl@aFlJlSe|eDlIl?aAa;l\\\"\\\",2):f(\\\"\\\"{b9l@l>lFa<l:l8lHa6l9a|e7"));
$write("%s",("lxb8a+e-a1bLf8aEfrl8arb|eidgi/l/l+l3a;ihi\\\"\\\",2):f(\\\"\\\"}l-fiikl=h7f6b-a+czbxbubHaqb6aqb4i5i3i5aqb-g-aff1bzb.b6fnbxbliThHgFghgHfkhxhckyjak?a=a;i;d*h3kziJjdh/ktcBa:i|b|bvbCihc=fUjbkGjBa?a:i6e\\\"\\\",2):f(\\\"\\\"}hrbMj?aKjTjwiHjDa?aEj2b3b6iBf+c:g-a8f-b2jCa3aKa\\\"\\\",2):f(\\\"\\\"{b;atgwbccIa3b1boj,b|b0adhyhdh\\\"\\\",2):f(\\\"\\\"{jSjwjCa:i.bci?a@izj>i<i@a:iyb3bCjyh3h?iwhxjBa>a:iPctihghgsbubwbTh-a3j1j:a;b.j1b0b-b3aAa3a7b-aTh.a:b:b,byhlhyiPaVh=i@a3a\\\"\\\",2):f(\\\"\\\"}hwb+b-aPccj/b8b1bPcxb;aBf-b;gZaWf|b.b5b-aUi-i3bDfvb|b6g6iWfMf3bgf;a<b:b3b-a8b6g,bxb2b2btb;ayhFhxiFh3a>a3a5anb-a4i/b3b4b.bHa8byb2bsgtbDfxb5b+bGgyhwhUhHhlh?g8f6fHapipiFaGaSh|fld4aogfi/ach4a-aMfKfMaFa=aFh-bHh3h2hGa+bJd@h9a/b5a|fCcyg-bPaBaob3h6aKaMa9aMaIa5axb3b.b4b0bxb+htbLfyhRfwhGaMb5g2bzb;azb-b7fccJa7b?a?achlhCdYaOaVafbVa"));
$write("%s",("ibNa=adhdh?a;aAgVaNaUaogchRfvbpbEa*c7bDaAaBaCa>anbJdubSczb=fIc?gyfwfuf2bsfNd3bHa?e-a-fGf:aIa+ctb,b:avbldub4bcb-btggcqgHaebdbJaGagfef8a1bxbwbtbxbUaac|b3bKffb/aRfggtbxc?f?a1aRf-a6a5bOf>azd:a,cNaOfwb.b;b>aHfob,c:a-a.b\\\"\\\",2):f(\\\"\\\"{bvbxb5a1aob,fCe2b-a:b1dtbHa6a/c2b/a:f-f;d+c1b/b3dMd-aDdBd@dmf/aob5a.d,d*d-b4b7eSc;axb+b.bbcZb0cbfJasdHa/aed+e0cGb/d,btb-b4aWbudpcgdLc=chchd6areOapc0cNb/a;bje/eGaHb5dedOb.a8aNd8aLdLa=a>aIaOaJapb6a+e5azb+cdcfbhc;aOaFdYd6aHaCa@aIaQd8aHa=a.cIbCbMd\\\"\\\",2):f(\\\"\\\"{cycvcocRapcXbocTa;b;bpbgbYdJaGbRanbQaJagbnbcb>dqc5dpbebnbOa8a0c4aJaTa5a+btb5bxbJaQa,c*cRa5a1bzc6aedMa0c3bldjd;aeded8ard5a6a5aedxb/btbvb2bxb,c1b4b3bxb1b0cocPa8aNapcMagdUc3b|b+b/b2b4arcFbnc4a=a?axbtc4aSbJcPbKckcic+bZb3b-bzcXbqcFb5aMa/ancvc+b+b|byb4a9cVbNa5aRb7cFbnbFbMapb2c.aMaFb."));
$write("%s",("a4a5aJaOa-a-b|b-aeb5aicybHa<b/akc>a>aXb6aOb/a8a6a/apb4a1b.b3bvb4b1b3b2b-b.bvb4anb/aJaPa5a8a4a6apbEb5a5aBb,b9a4apbpbnb8anb4aGa=a:bJacb!5R1ca616R.ba~[2xha=s,y=z,54[54%.4[e6&yay,]99999[gnirtS wen=][c n3aea\\\"\\\",2):f(\\\"\\\"{)v]y3b&a(niam diov citats cilbup\\\"\\\",2):f(\\\"\\\"{RQ ssalc~5[~5qfa cdlnl3c/a;maertStnirP/oi/avajL tuo/metsyS/gnal/avajq5bdateg@3doa2 kcats timil.v3dga]; V);U5aC3ecaL[f6aa6hha dohtem?3e;4nga repus&3ecaRQ@3cgassalc.@6[@6ioa(=:s;0=:c=:i;)$5ajaerudecorp34[34eqa(tnirp.biL.oken\\\"\\\",2):f(\\\"\\\"{24bianoitcnufc:[83\\\"\\\",2):f(\\\"\\\"{martStup=niam^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4)"));
$write("%s",(":f(\\\"\\\"'>3(ba7U3vJ4vba7I4.da,43?4[fa(f;)5/6/#6[#6[#6[#6moa(etirw.z;)tuo.-@aba(q?b~auptuOPIZG.piz.litu.avaj wen=z|5[a7[a7;ca34A4.l41ba0j4[w5ada283m4[x5[j4fea1982m4.batv9[V:[?4:da12927[=8[V:[x5[x5vca04V:/5aR0Z0Z/512152353/2/2166263=4/3141726??:1518191:1/I9[.;[?4:da063.G/r9[/;[x5[j4Fda66957/da*6 .C[Z:[?4;da348Z:[A8[Z:[x5[57wca8457/ea1312aC[a;[?4<da423VF/C8[a;[x5[j4Fda200a;/YB[W:[YJ<ba1OV0>8[W:[x5[YJGca15XB/fa41310\\\"\\\",2):f(\\\"\\\"{9[[:[.[;ca92B8[B8[[:[x5[x5wv5/qa;t:\\\"\\\",2):f(\\\"\\\"}%%%%\\\"\\\",2):f(\\\"\\\"}fi\\\"\\\",2):f(\\\"\\\"}*-84OH2ca7786[86[Q8[x5[QPwba9R@/(a]i[\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"}+17\\\"\\\",2):f(\\\"\\\"{<84.;i:-i602\\\"\\\",2):f(\\\"\\\"{;i:911\\\"\\\",2):f(\\\"\\\"{;j:6323?[tA[?4:da550d9/xa(tnirP.tmf\\\"\\\",2):f(\\\"\\\"{)(niam cnuf;V4[;6[;6;ba93;[><[j4gca69mO/datmfY6[>8[5R;ca5847[?8[V:g"));
$write("%s",("ca02?80saropmi;niam egakcapo7[O8[?4;L[1ga(tnirp[A[+6[?4;ca36(I/|<[j47da444l4.ba-W6[<8[i<[A?njanirp tesnw41ca21T9/la1 etalpmet.f6[F7[)L<l;/ga(ntnir|D[*6[?4;ca93SG/baf)6[)6[?4?ca11EG0$a,s(llAetirW;)(resUtxeTtuptuO=:sc5[C6[?4;8=/#BaC4[(6[(6[v3kdaS C&6[&6[*D<3=/ca&(?4[$6[G9[v3kba r=[)6[)6[r=[&6[r=[83)iaRQ margoP9[-6[-6[P9phaD : ; RW9[-6[-6[v3mba^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'>4[#6[#6[#6[#6[#6[#6\\\"\\\",2):f(\\\"\\\"}i=[$6[$6[v3lqa. EPYT B C : ; A36[36[36[y=[#6[#6[#6[#6[?4[#63ka)*,*(ETIRWs=[.6[.6[G@nhaA B : ;,6[,6[,6[v3lba [2cF4[+6[+6[T9oia: ^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\"));
$write("%s",("\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"' ohceI4[.6[?4[73kpastup\\\"\\\",2):f(\\\"\\\"{)(niam tniL4[164ca01?4[?43ea%%%%@4[%6[?4[%6[%6[?4[73\\\"\\\",2):f(\\\"\\\"}paparwyyon noitpo26[M45<4[<4[<4[<4[jD@hanftnirpD4[fa(f;)3D4/kaetirwf:oinu41ba2u4.ja>-)_(niamt4[Q8[<4fWP0gacnirp(C4-ia(stup.OIK4/rKajaM diov\\\"\\\",2):f(\\\"\\\"};)B3(ca11g62oatnirP)--n;n;)sn3a<a(rof\\\"\\\",2):f(\\\"\\\"{)n tni,s tsnoc gnirtS(f diov\\\"\\\",2):f(\\\"\\\"{noitacilppA:RQ ssalc[k4rga@(tnir>MblaM dohtem06x*3cl;abNcuadiov;oidts.dts tropmtNnra1(f\\\"\\\",2):f(\\\"\\\"{#(rtStup=niam&3kkaenil-etirwb8dva(,^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\""));
$write("%s",("\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'s%^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'(gol.elosnoc;)^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'73g\\\"\\\",2):f(\\\"\\\"}a^129^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",12"));
$write("%s",("1):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"' nioj.)1+n(yarrA>-)n(=fI3cva^31^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",2):f(\\\"\\\"}54,1\\\"\\\",2):f(\\\"\\\"{.^127^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"# qes-er(K7c.4cba^31^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"p3lg3fw3hla1% ecalper.j4dea^128^gXc/arts(# pam(]YALPSID^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^127^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\"));
$write("%s",("\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\".NOISIVID ERUDECORPA3cma.RQ .DI-MARGv3g53d|bNOITACIFITNEDI^127^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"[tac-yzal(s[qesod(^63^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"))System.Console.Write($^63^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"Put caffeine \\\"\\\",2):f(\\\"\\\"{(int)c\\\"\\\",2):f(\\\"\\\"} into the mixing bowl.^64^n^63^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");M3pva^63^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"Liquify contents ofE3oeaPour^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\""));
$write("%s",("\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'3w^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'4e\\\"\\\",2):f(\\\"\\\"{abaking dish.^64^n^64^nServes 164cma\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}^31^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");\\\"\\\",2):f(\\\"\\\"}/****/e3a^15^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"),s[999999],*q=s;int main()\\\"\\\",2):f(\\\"\\\"{int n,m;for(;*p;)\\\"\\\",2):f(\\\"\\\"{n=(*p-5)%92+(p[1]-5)%92*87;p+=2;"));
$write("%s",("if(n>3999)for(m=(*p++-5)%92+6;m--;q++)*q=q[4000-n];else for(;n--;)*q++=*p++;\\\"\\\",2):f(\\\"\\\"}puts(s);return 0;\\\"\\\",2):f(\\\"\\\"}^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"))\\\"\\\",2):f(\\\"\\\"{s+=^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"00g,^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";for(m=1;m<256;m*=2)s+=^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"00g,4,:^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"+(c/m%2>0?^7^\\\"\\\",116):f(\\\"\\\"\\\\\\\"\\\"),\\\\n(\\\\\\\"\\\"\\\"\\\",5):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"4+^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\"));
$write("%s",("\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\":^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")+^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\",^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";f(s);s=^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"4,:,^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";\\\"\\\",2):f(\\\"\\\"}f(s+s);for(c:Base64.getDecoder().decode(^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"kaAREREX/I0ALn3n5ef6l/Pz8+fnz58/B"));
$write("%s",("Of5/7/hEX/OZzM5mCX/OczmZzBPn5+X/OczMznBL/nM5mZzBPu++fPPOc5zngnnOZzOZgnBMGAW7A==^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"))\\\"\\\",2):f(\\\"\\\"{c=c<0?256+c:c;for(i=0;i++<3;c/=8)f(c%8);f(^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"8*+8*+,^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");\\\"\\\",2):f(\\\"\\\"}f(^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"@^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");^1^\\\"\\\",4):f(\\\"\\\"'|sed -e^1^\\\"\\\",4):f(\\\"\\\"'s/^16^/^32^/g^1^\\\"\\\",4):f(\\\"\\\"' -e^1^\\\"\\\",4):f(\\\"\\\"'s/^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\","));
$write("%s",("9):f(\\\"\\\"\\\\\\\"\\\"/^16^q/g^1^\\\"\\\",4):f(\\\"\\\"' -e^1^\\\"\\\",4):f(\\\"\\\"'s/.*/print ^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^8^nquit/^1^\\\"\\\",4):f(\\\"\\\"'^3^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")\\\"\\\",2):f(\\\"\\\"}^1^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")\\\"\\\",4):f(\\\"\\\"');\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\").split(\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",128):f(\\\"\\\"^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");for(int i=1;i"));
$write("%s",("<a.length;a[0]+=a[i+1],i+=2)\\\"\\\",2):f(\\\"\\\"{a[0]+=\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",185):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\".repeat(Integer.parseInt(a[i]));\\\"\\\",2):f(\\\"\\\"}System.out.print(a[0]);\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");\\\"\\\",2):f(\\\"\\\"}\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";FORiTO UPBtDO INTn:=ABSt[i];print(REPR(50+n%64)+c+REPR(50+n%8MOD8)+c+REPR(50+nMOD8)+b+\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"J\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"+a)OD\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans c 0\\\"\\\",9):f(\\\"\\\""));
$write("%s",("\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"do\\\"\\\",2):f(\\\"\\\"{D(Integer(S:get c))\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 35 39\\\"\\\",2):f(\\\"\\\"}(<(c:++)(S:length))\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 24 149\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");end;\\\"\\\",1):f(\\\"\\\"\\\\\\\"\\\")\\\"\\\",1):f(\\\"\\\"nsys.exit 0'}\\\\\\\"\\\")\\\"\\\",0)]]></xsl:template></xsl:stylesheet>\\\":s=\\\"   \\\":For i=0To 7:s &=Chr(32-(Asc(c)>>7-i And 1)*23):Next:System.Console.Write(s &n &Chr(9)&n &\\\"  \\\"):Next:System.Console.Write(n &n &n):End Sub:End Module\")\nput=s\nprint\nqa!"));
end endmodule