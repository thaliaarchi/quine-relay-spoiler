module QR;initial begin $write("%s",("Module QR:Sub Main():Dim s,n,i,c As Object:n=Chr(10):For Each c in\"<?xml version='1.0'?><?xml-stylesheet type='text/xsl'href='QR.xslt'?><xsl:stylesheet version='1.0' xmlns:xsl='http://www.w3.org/1999/XSL/Transform'><xsl:output method='text'/><xsl:template match='/'><![CDATA[write,format=\"\"%s%s%s\"\",\"& VbLf &\"(\"\"\\\\write{-}{txt}{(\\\"\"with Ada.Text_Io;procedure qr is begin Ada.Text_Io.Put_Line(\\\\\\\\\\\"\"print\\\\\\\\\\\"\"\\\\\\\\\\\"\"STRINGz:=REPR226+REPR153,a:=z+REPR166,b:=a+\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"2\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"+z+REPR160,c:=b+\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"8\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"+z+REPR165,t:=\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"write('implement main0()=print(\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"BEGIN\\\\{s=(\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"#include<stdio.h>\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\nchar*p=(\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"Ra#include<iostream>!nint main()\\\\{std::cout<<(!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"class Program\\\\{public static void M83apbSystem.Console.Write(!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"let f(c :Int):Latin1=if c=127then!!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"!!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"else(string_of c@!!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\" g caffeine !!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"@$3kEa!!!!n!!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\")@f(c+1)in print(!!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"Quine Relay Coffee.!!!!n!!!!nIngredientsq3aha!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"@f 10U3cgaMethodz3c#a);let g(String ->[])!!!!n[c;t]->w4edaPutY4spa(int_of_char c)05auainto the mixing bowl|4ejag t!!!!n|_ k4gtaLiquify contents ofE3oeaPour\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'3w\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'4elabaking dishv6biaServes 164doain g(!!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\")))s!![2aca!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\" [2bo3cparts(nltnirp(])]v3cja.NUR POTSp3cx3dp3jba!!M3dp3df4fda[))j3ci3e,3cp3l[2kga\\\\};)06xu3kgaqp]\\\\}\\\\};@3\\\\}ga)1(f\\\\{#+3~ba3+3&ga7(f\\\\{#.,3~ba5&4\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'ga13(f\\\\{#+3O97l,3tkaD ; EYB RC73(da,43.3\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'daDNEZ3Sda. Ab5VeaPOTSc5Wb5TmaRQ margorp dS@aj4ObaSj5UV3Lca36V3Vba&P5MX3agaS POOLi;Vea\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'&,)i;Uga. TNUOf5Tfa(rahco7Nh5cgaB OD 0l;Uca&,t9Rca)At:Vo:UiaEUNITNOC0Kaca01r8Uk8Vn7OyBceaRC .b4Ska,1=I 01 OD4FWcaPUc4Tx;Rva;TIUQ;)s(maertSesolC;5Qmr4<la721(f\\\\{#n\\\\})8i3ag4Mda531w6&ka(f\\\\{#(tnirPwS$Y4"));
$write("%s",("Sia115(f\\\\{#\\\\}Y3Mla3201(f\\\\{#mif/5$h8*da402i8cj3bi8Mqa904(f\\\\{#;)\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'\\\\})8225w8Tta75111(f\\\\{#\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\',\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'&\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'(rt.\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'&:Nba5x5a\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\':Qba4RW,w7,eaq\\\\})6j3bh4Tg5Mda728\\\\}:\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'f7-ca96/>aca\\\\}\\\\}0<Nb6Uj8[ha!!!!\\\\})785:BUea9052i6Yea&dnel8[l8Tba3eJ\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'$?.ca67gKQh6[$a\\\\{#&&&PUEVIGESAELPn&&&&1,TUODAERs3amIMca70#7Uba5pIb;>[FC[wLLca48:?Uea3522/9b~a(etirw;\\\\};u=:c;))652%%)u-c((||~6[*8[4;Kba9yLUea5063U>[ea&#-<k8[Y3Fca93WCVda757l9[t;[ia\\\\{#&&&||iy=Nca38GW(=?.ba1a4a\\\\{>[n8[9XMba88XVca23\\\\{>chaBUS1,ODh6[p8Qca82*N(FW/+O[$>VVHbma)3/4%%i(&&&&HT[LXHca632?Uea92713>[\\\\}8[fa\\\\{#&&&/TRda701&PUda989CC[o8Vca32X3(MF.ba7o9[-TdNa2=:/t;2%%t+2*u=:u\\\\{od7 ot0 yreve;i-=:u;1=:+i\\\\{od))1(e"));
$write("%s",("vom(dro=:t elihw?s;)s*hU[c9Sda254$?Uda546q<\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'i6[iU1GI[k=Kba4u@Vca35u@a*D[wXRba5u@VFMaHJfg6[*D[h4Jda197$?Vda031&>[nb&n&&&&dohtem dne.n&&&&nrutern&&&&V);gnirtS/gnal/avajL(nltnirp/maertStnirP/oi/avaj lautrivekovnin&&&&u9[u9Rba56?Vca146?ai6[u9Qib&&&&\\\\}\\\\}\\\\}\\\\};0=q;)]q[c=z(tnirp.tuo.metsyS;)0(tArahc.y+z=]++n[c;y:]q[c?n<q=y\\\\{)0>2%%++i(fi;48%%)31-)i:3c&as(+87*q=q\\\\{);87261<i;(rof;n)rahc(+55Mca74I[Uda126?:[jF[?ZPca42?ZVda481?:f[2cm6[u8[/MKca69.MUba314aT?[[2doa=]n[c);621<n++K>aqa0=q,0=n,0=i tni;<8[DJGca36R?Uca56=9[E;[<8mgc6a2b9a392a4a5azb-e;axboCbd,I6aDdehLa4abdZcFEN24aJaJaeh-ar7-pA+HaPdTbpbZb>aCR51>,/x+bIg/x\\\\}bJaMa\\\\}bJaPaIgG-JaJacdJaJaTaJa8bW,;ad<TaKad<Ta5HIgPSxSSamE9bKad<3JTad<d<Ta8bmE0qJaLaJad<8bmEh4cma8bmE4bmE:b/x&4cga\\\\}bJaHa\\\\{3aca0qk3a@b"));
$write("%s",("JaQae1;a8b>P:aUa:aW,CbSiNcie-awbHcFcCcAc/aZg|bKI9cYb4cYj0c|bKa,c=auc@aEa0c*c3b|c5a?bycc4?aYBJa|bieVbpbTb;g4dWdpbZbHakcHapb6a6a9c\\\\{e=a-a-kOc3b9d6a6ao3ada|b9i3fra*e7apb>z7e5e3e1e9m3d:aShTc1bS2Bgpg+bWium7a>z5a2bOhMa-kOcufvbJa>a2a:b6a5a-bHy3bia3fa<gd6a53khb9d<dvbgdTd=a=aMdXe2=-aRa2=kbUa92af>eMeaf=g7bmfeh9f=gIcGcSgLhggQhmfhdqg4b-boi9a4a@i@i4amf/b9d;adJQoa(f\\\\{#gfbiVj;gt2F6a44a>:c-a9abj=g,l2amfmq=gaf4k|i4a4jLhggJhJ74b0b9fy3cia@i9fpbYeo3e*baj<bSg-i9d=gciefDd?lJ7g,Gawfnd+b-VSV;a,bWiT>fbpbYeA7R?5qhrnb?fXfAY5g/fufvbliBiWh4iUhMgEaElGgEhChdg9a7bed/f5b<6-bCh3a=a9a7b|Qs3g53ecaCh53kG3a33iia,b9a7bXcs3e\\\\{aTh\\\\{8xi9a7b+;/f5b.btH8h1gai53ak3a\\\\{a/f+b/e-egfCh3asbDhEa3a9f=gq5eiahhDhCacgs3gcash26coaggBi2iAhyg9f=aC7eG3ica3eC3i5agi;i=gygwf:bSg-i:\\\\{392a2avnmfphtj7gHc9f=g@a3c=gp"));
$write("%s",("br:a1a;gJaJaubzcmfKf=anb?f<gqhyb<hmf,bJa=g7b5aSg-iG3c?3esa9a9b9a,hagqh/f=g>aq3aca5eq3c1a@auc|b9a0b9a@a>a7a=g@a>aIa|bmf:a9bJa0bagqhskW3c%a,h9aCaAaJa9bagqhYfJa6aSgtimf,b9fo5gyauiQhBv/f1eSgRdpbYevn/fvnQ3avasgmfbqne/fvnoUbb/fvn/w=bw3glavnnbggJhle/O;b4a;g9a8b9a7bmfMaJayb>aB-dDJa|b/fLc9fygwgJaj\\\\{dDJa-s3bda=g=DEMxa52(f\\\\{#(ntnirpn\\\\})821(f\\\\{#~>#n40+ag@a>a<a2bmfMm>d:axiJaubmfqe>djn4b-bJa32>fkaggBiyiwi3aL>e2:eoa1i/iwbHcDhXj/i\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'?b;ak6i?i=i;i;awbHc=gvn?.peBjyj\\\\}lEk\\\\}iCkKlhj5jOl1l-a\\\\}iQlslTy3d&j*jk:ioRaubzWR\\\\{wq3A1A/ABaEa<oBaEa\\\\}bxOImcp\\\\{AkT>zSaTaGaLqz/56Oa,|ln,be-6IibSa:u<u0n|obul1om,0>a\\\\}G+b0*9b7b\\\\{8DmO,=aBak:n=hYK/0*9bEGibCaMUibE-o|,u2bkTDK\\\\}G5ujb5b<9HJ,\\\\{e>SaZaC<0bUS7b7;Ea/L3Mj7W*ib7zB4YamboeHv?.7m,b04mb3n.b3oAO@aBK5bmbhmmrY/UaXa\\\\{LB5f"));
$write("%s",("uzbc\\\\{eb-bnv+ryDu,WavbwvA\\\\}/HZs9UEwsNZUF?9gZavxZ/q,FDe8YaPx-|QDZkIm.b?3zbMt-bvG+Iyn:5@aAnk--u/JSotmYag3+kzWE3W*Na3bu|Pa<Dw|SCyMTQH|b+5mUa<WEa9g/bsrQOzbgZH5uS5bibcXfb8<Ya,?xFFuCats\\\\}-PpQz,S\\\\}mVa50,bIcA\\\\}ab\\\\}Nep=uAz0bx+l-b|.tqu=B6/bbA+Qqr7BpZaznH;XybbrCtsNaj1J2BavneU===JbugoDxI\\\\{\\\\}/RaxWUCcp*ohb+tO|\\\\{5TteO9U1bFnLScnOa+48sQadb9u5GOaAuzpxOKnmQs0-|6>Waus>xubGAjFDaVa9gtbEat3N-NHEal1om5bR=*oavEa5b;G/?BaEG=BZQ\\\\}?lbim5S.bx?imu?ldr?,bMUAOTa9>=CB/<a,bTunt71Sa,bcnmbjbB63bY>JSV>Sa,bS>EadEP>M<H\\\\{jbR1Ra@amblbXzwfCFD>m=gZVqom.nLFW.m?|mOW|bmnP0ibvz|m-yV\\\\{lFhHAvywsD3zp+lb?.Bau*1b-b@yT3gmkslGUmDa=c0*c3c\\\\{e0?>L|c,b@y2=EaRcdXb>4rTa3=An/t2=Ea>VgZmmA,41Eav=fbEttx@y\\\\{mF=3toVEG@=<=om6b41Ea46\\\\{>lbtp;vZa0=3zV0IUEa6bR?@y<6dpI:Fw41Yls=lbzb\\\\{>j7n=cbl=;vzbUMg=;vwt@,B8fbd"));
$write("%s",("b+bAa\\\\},+bAaxZibCaYa,uFmfxPuMUTanDSa,b@,av\\\\}GE-Naj-0*\\\\{d0*YQAaG<d/D<EJdb+bh0\\\\}b38g3xZ,qFaFywf?awv,bL1UVi\\\\{x:*G:5Vo;nftorstN-9n,<\\\\{8dL,bdb+moustj;E|eLib7b:5xpHYywDa0b<a>a;G2e0bGoTa3vb,DapnwfDzTaXa.bnnoOpnwfR=9nH62s:51iR=<aWrv\\\\}Tr\\\\}3cTd\\\\}/SaZ/nn<n77X\\\\{z|s4hbRa12pKW,DmA965J7:yoO/;xb6@db1C2MjH3nc|\\\\{nfb?ab4fb4S2b\\\\{/7bPab+g;abysP7S5V2abUZfb,s5-2ALSy/1b*by/CaOa?av=fbYz0u0?v8N-d8Fa+\\\\{,\\\\{RaABmysSqs7bo5z.xw<a=aTaAICOCaKnQ@E6ibhmvbmQUts+Xz\\\\{bnK-bd@D-,o,W3e;nCe,W3ePZb+hbRadxQvqrg\\\\{Br0iO=z|/tB4KPizZV;/kTF,m+<,3b+F>xW\\\\}Szbu2M8biR.twbjTTz:p1bV:>03fgur|9b1bkbzPkfiN4bor2sd\\\\}Aq|<m,4b9bIxgby2K?GTQ3E5fZatbvbFajuwfcXYauo9tCKgIJkh1CHybE,xQ>aoL-bhb4x|J?.Fax?gd\\\\{mk85YGZ:qT0|-GascN<b@5-Va5m3mXw.n\\\\}qsrXHn/u>-|>r/b-qJ|DaPCioY/?ron+FfdPuv4uw.povg75Gan+G\\\\}Gfd7DUA"));
$write("%s",("B\\\\{/oUvJY9b7bQrrohbrCuw4.Oa?air/r2b0pgbj7i8TZbb/pP94t5fRai8ab|*Yarxltcb-X,EYcduA*>9@aybgCh0G2/b1o,btNEwB\\\\{9bTeubP4P9b|?z-pA>X1nQYH-7VzbbebabjbGaEzZ<y-hJ9bXcauKqO=GmVe-21H0bRBNa?.zbioQ3oBZaVETEEa<Ga+DafbMntqgdSf>Bk>Hcroz/Va\\\\{>4.6C5bib2bfvU-h1:vZadTzbh1:vDaZa>a2sG+Fa\\\\{4ZM3qUat5x*Tr>a2scp\\\\{|1vQFRaS\\\\{\\\\}w6bRaHc?aKOpGAOxZJ9cpmE4bH/aB+4U\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'tnirpWMNga02(f\\\\{#LZQba4a4aja wohsn\\\\})8o3bo5Mqa904(f\\\\{#;)\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'\\\\})6307|5T>g9439(f\\\\{#\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\',\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'&\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'(rt.\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'=kb6J41i*C=2B\\\\}mYM1vzDYQI-;pd+Lzl1gbmbQmHv\\\\}wx*ntybPah9ubV+asauu1ZaGtv*/:b/sNxQKnB89QM4t.\\\\}n2b*xGx7sNp0YGx.bd@9Q1b\\\\{6qn0no7PaUaGr*b<IFajwlb1m/bjyJCyO<>+q3b+I/b1bf9\\\\{bC@o=?ayb1pMuM\\\\{-uv\\\\{gbFad0Tt8tR\\\\{@n?PTaG4Ppny?p@a.X9yjbPO0bQDC"));
$write("%s",("<8+evcbuI4@sss|Y4Ta4E\\\\}74@@p>zfpHrz/-CA@QD|J/N|p9|Va?a,ShHXaRt?<x\\\\{U6<a5bBaWao/>vhb6enywlKRnvY/H.QR7blblbp*R\\\\{l>Xzcyu;KnxP6b*Gb9EoLEbubbMH|Q79\\\\{bx|W,V8as-bWaf-A@C\\\\};17bwbKqIoA@*Mt/ymE1BaaBP@jbBaed<u?rkuYQ1t=LBy0C77z5\\\\{bbfB/15x|Zabb34eb-bpyeb4e\\\\}b3=Ra|bF2ZQ8b.HV\\\\{5bUaZc=I<hVenNd/<xp56PIF@qltKqR4ov0bGa8L-FcbVf.HkbPw\\\\}DDzNOavz;//ZQ0bL?kbPwwf/7\\\\}J\\\\}gaL*Xb4a.kgqhbzp?*V2UiPzj;lbRa\\\\}bXM7pMfabu4\\\\{>oSow7zQx/b|pNa\\\\{dU6*b.Vwf/72WTa?v4+*nKtbAkbI:Wp+Ndm<Ayst.rZ16I-HJ\\\\{.n54bou<a*ye=6988Ir\\\\{*W,.EBadDGa\\\\}MWNMpsN.b6b/UmJcbY-Ba4bQFFuHJ47ptibFaPC*9|t?rq:6oNOF,ls<akUO.mBjbp=*rCVNakbyb<uoP4bD>OafsRve9@\\\\{AqWaq:fpj=.1NaS+V2|\\\\{|tN<y2-oE,ubQ+,WBY,b.b8.9sXvzAiE9s;+=9fbq:+bsxPa7rNaKIQD|buV4-e8K|Zagix6.z2S|Qp6b/Y1*pYa8b>aoPqmNa,bf*QaO:=awfCRg*oi9,23E3C6UvO0RRGaB,o"));
$write("%s",("4.b1v>,-qirhbNXbwEhHtE|5b+49171+W;077db6evX0mqdirly5btU;M+X\\\\}mD1kSioPwP@<|?a>MsyH3.Jwb-:*ozbCt,0y4D4Uao/w,HTVasW<Nvwfm,bwU0P.bCt;ISG5bc7uXCmFa5bwt:s6ohMQaRa6brD+kp\\\\{o4\\\\},9373S*e76CcbQa*bwbw0jt8\\\\{vb@+?8\\\\{bbbhb;M?ap*?7qKNaMtA/:|1pNpG9?<5b41jwDa5x0m?E/b8B=;5W6b3W/PG|z;LVSaSV.p+41pW,*bJ3C=4V6>*Owb|OebaMqD/bp\\\\{wfNHSnOptqJ/6/*G*D=1n,.UpOUas<y4\\\\}bt|nKeb?aTNcteb.MnyPaV\\\\}3NsHCqu;NFcbp\\\\{+rzb/w9q7qWr2-2bE3L5q49blbUF<vib\\\\}gNFYa6bzbL5zbP<pUEJtb4G.bhwbbd0x5WSCaVH?5pVC=SKEgbb?a+RY|N\\\\}cbJwyb\\\\}b7:-C@L?yy@>wv,5vx5k-qo:t-bSuwbBaImstX4Eg45PC*GF@jbDaYa-bqEB+GQc1(f\\\\{#afrzdSu\\\\{b+w+v\\\\{,CRhMXFR:?<:t>L+,Oa13U6b4bfNabvA?qv2bZa6bYoSfmzi1Na,.op4@Aw9oPn0iin-beCvGjw*b.bvpty-b+zFmopF?kl;\\\\{jy9\\\\{Y?Bv2@Bv+z\\\\}bgAUo*wjbi\\\\{tKy,8b*RjxHJ>dtHQw;Gwb8bdbyq;IdbR;aq\\\\{,Tab*79Zrm:6"));
$write("%s",("Bq\"\"),\"& VbLf &\"(\"\"sr?l7NNynoLMFk-Va-+3bQ\\\\{CP,p3+y/O2D.p,dbV\\\\{h1FaaTezJoA;.13Q.b4b\\\\{J>a7SkbYa23l6qD9bQaWa2o\\\\{6S0Cue+6b+bL-/twK>CEh32PawfW\\\\}DaCa/+Tae=H5TvZQibQAeb\\\\{3@,JGA+IoL\\\\{<>9bzbFye-DaGaz?NaHvPa|b-Q9b0GFa8bX+ImA*BHE@9bs4SaPa?vmbC.ZapK4RRa7bqyUa4p?.?\\\\}1>t/r/6o98+>wz8u3q16qRfb/NeRPw+o4RrATadtY95bVawzWapCOaa5WN6x\\\\{R>a3bP3@anvNa8ueb4LasWc|ERa9g//uRMpAaWambg>mblmNqV94bwfmEZaPM|,N.R.qRUa7b9H8b1nmbzbU6TaXsUaa,qIQaX+D.B.Rac7s+abX>,b+bo@PO/sJ+VaHJ|,J2w\\\\{?p\\\\}04tj7Kmau4@wu+-YHinu;ju-QZ/j;UaD4RoSatF7bmbDwjbJog4x.<aBGXMiqbxCatbt330u*=Kxbv;8ojt+bR:?.Yaw88bUm+-FD1b7bBaxBenIgw4Mf6b?adD=aEIRcKPrr?ClCCKx728axJ+AarxDwWad1Fao@Da=as+aPF\\\\}.oR1NpSaU6AaK+SaUaAam*NaSk,?17H1=a6b=-.1\\\\{A3e*5/binvbwmgbuPrOIvxPWav,6b8qn>WzhCWa,p+bTvwfQa3>vb7851UOx\\\\{J?-1yD9t8*g7Ra=akO9"));
$write("%s",("b|458RaD\\\\}2@epybDa8./bf\\\\{eb5b7busU=@**bA*M9Ua2-wbv-Sx\\\\{b+ou6gmJ0g9d+XakOlr:?aqa;CKT:l7\\\\}bf\\\\{GfwbG:J?0b\\\\{@?.NaubFET1n>mb/7\\\\{b*b?aDa<FO*9=TadKOw=,?|n2cb6oi8:qqrdqbqE4Zau372FaR2-|fNibwv4-C@8p>u15+w,b8qAanzl*9y\\\\{5fdiv6eubdNAa1b+=E3S;YqGasq6xGaU2QrHqmb46zzRa,bn/ibl21b13p\\\\{;rwfP?vuVn3bWBNmmDDx7bkba-=:\\\\}+tb1mKI*pG4eb:rtbVn.bhbUazuCeztcpn51>f*5bK/ybt4p==:pCSa4b>\\\\}\\\\}Fs4tKaw\\\\{p-|Hx1p+Mir63,bmbQay,cb\\\\{3duGrwbzbXvwdsy?.bb4I2bwf1bO3qDcdzbvJ4Lw*VaXmXrOLML|,h9xx73ibabqzX\\\\{+bv.AzGn=;>L<h2bO2abfI-bC<<q;5db+4r5y@d=1bExFnw|WCXFeb3bP<Vf\\\\{>.nXF\\\\{dLpWBYaMF@+U15K;zNatK@,g\\\\}Aafb0bH61nCaRq|r5xC6q/9b*:cbCej1KG0wzyjt/rywf*cqJsSafb1,g7L.hL-eCjyKwK7b<albvKlb<mdtSKt4Sk4b,|7b?s:KO\\\\{50By/.dpQa763KjI=*a<0v>aablb50Z/Ra4-ub?.Qa3brKemQ,NaCamzSa3*fx+nW:k2D-Xllm3*Va,ype<mSa"));
$write("%s",("ubbbl1vbjb+nZaib=aHtebaKg9zbexl-UaCwa<,|5bg=,y+bus-p>mPwN=n,Mq3*2>.b>a@w<6506/Dvr:6oFadfrvfbUC;o1p\\\\}n=4.bkD2bYmmyRabbr98\\\\{wb4vN5?ao;Ua*bZayb73@6I:@mRakbUn@a2byb>\\\\{lm-b-bv7\\\\}AL?A9*bu*\\\\}bd\\\\}.4J.TatFjuCawtw\\\\{L5|b/rKI.eIgqo\\\\}wsIUa<a3GW\\\\}OHMHmC|\\\\{*b2b3\\\\{C?ZAsyZFeb*bexh\\\\{?.SaPxJqabxbhbf=5b+oRaFm\\\\}b-bK5+@Ixab6Co02BGah8ao6:kpT34E4=8b=:N2<aw\\\\{bb6rFDz.K\\\\{@ycwE4b|mb*\\\\{rxZnEa=pMt2bd,N9h0wbR9mbybPCMA0A+@W\\\\}-biw/bYaV,P\\\\}K?d8\\\\}bAax.EsguSa7wybT6b/@wRa6/1>-zRa4p|c8bTa9<Q+ZaO?s<lbfbye>zUohbmbn/PCN.ZaVuParu,bwfKnLwu6=tcbooGaa/J,Fa|DjbXrKvO/ybXD\\\\{bjq.@<a.?@,Ct\\\\{,S5-b?teqcqU1;n85i1g1<aZa-qE@5nvb?.ZaDx-owb52b@52\\\\},jbe-as-7FEt,Zav.FaB\\\\{42ebrBP@fr7fczYadblCvb,pQE-f>r>albS5>as1-7lbF47b?Ejb8q.@bxdEKqT-d8K55bJ\\\\{T:Pak.gb<dD>e9A\\\\}:pIFtb*bD>fbjbWa7;J;RaLfDr6bh"));
$write("%s",("\\\\}?a\\\\}DAa8FBrPar5<d*bv.o|XauFCa4bEa,FH6hbj1=\\\\}x9EalbabgbT<;r2bMpzp9Dabo\\\\{<xA|Ya>av=g*J2jFh\\\\}ubcnnpYaVuyb+1?728>a\\\\}+o@:oo@6CKn?CTaWagbYaI\\\\{Fy4b/yT|-oA,QrXa?.d0ri-b@a9oW+t4PwLoYa,nY9JARt0b*yv\\\\}b+\\\\{bRD2b-sApvu>azbvb*Dy\\\\}O>ybaBTa.ow,<a4bnEbdxbgbIr+oym9zqepx+b*rEt1iQaJ?R5VfO3\\\\{bs2>a@zXvzbZaAB7bR;yb=;o\\\\{wbbnAr-2y8wfZ/J\\\\}-bL\\\\}h/gb-7\\\\}Ag\\\\{fbY9df2D>vwAvb=|hbCaAntb\\\\}bgbc=Y5b*W+nw<.b6=CA3CaGa+:ibS1pqXa;0@aA\\\\{LzlC5bU-<a-m69\\\\{bmbA\\\\{+b5*t/+>EtxpGavcvw+-=p5fd1Za46Mrmb\\\\{rNaKqQq7bRa1bZl.58v>=X\\\\}+b7bTvlwWsawfbDoJoxbEa>a*bwsJo5oTa\\\\{tmb?a=/9b>aYa*b,0>6yb6b9opiLwEa?<Fa+q82|bg7kbO1botbT=+bFfL4QaubPmSaYz>a6b-q|bwmH,ybYawf=awbUaGa/n2br5\\\\}bz/vui?JmzA<aD4W+6>H0U-0AXqV;,w?aOa\\\\{bjBC67bb4.z4bV\\\\}wv3tublt2vRavb6bCAOax*l,+zZlH8piDarxfbbb-b3@ubGaQ5C=ub23Bvl2uo5*"));
$write("%s",("wv.48.*zG;=,+oU,u?;mwtmb0b@/2bTnpuTaXvwAGaBcH;vptp/beb=a-bZ/v,Rak??.hb=;ByA2vz:q8qv;/bioog.b8o1bwbXa,0Qx7bk/abY1,Ah4P/e<C=Fae=/bDaV+Ua4bXaA\\\\{<aPabbAw,|jb.ze-bokb6eXajr/bubb4o<4b1bi\\\\}=9<wYpGeGa8zEam:/b0b2bEw-ukbirXzR967Ur6bybRa|\\\\{wfl10b@aa\\\\{Y/gbarIc7b1uTnRnyvO>Oa,bVaLt46wvWaA/\\\\}sZas||\\\\{wr9b.1abOa\\\\}bW<Pwb+9ginOvVnAa32X*Yr1|k/;|VogbH9WaYaTxjbk2,3dbpqP<vb9bA?Ig1bK?cb=ax|P\\\\}fbwbib<=wf-uQa0pe37bRugbxb?.+b1mJ:*p7mf\\\\{UfuoQ3Sn0bk/|3T3vb=,Xal:Dapquo9zw?b/.bNt71/b3nvb,bqrybw6hp@albUahb8bhbgb4828=,+=F-Batb@awzq+6/3b\\\\{b.z8bZodn0p7zUa9dUtc\\\\{Waoyvzn|ab3bTx>a4xt4wbwdjbV,;=xbbbG,PaF<B82bMttz@a@wlb@amerrR,b+bbx<db<wfb=pN\\\\}p=2|H=3bomdd5:<ajb5:6b\\\\{-4bVav,R:UaN+Z=|bX=*,x\\\\{X+,vRc*,ab1b2bQaC6-bEt8t?aSavbW.IrG;Sahb-qy0iovuYal:Ra82vn:\\\\{sndb6=F\\\\{K.6bR;kbxx0blbOaasP"));
$write("%s",("+R;LslbXakb6bQ+gbny3m<9grydRa.m!![2aba!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"g3b[2lpa\\\\})1(f\\\\{#(tnirP;)23&Z02b2uj=09xb>aPawdUae=|b+o8sUabbOaPafbydkbubfu+kZa2bk\\\\}wbEgFrp5Xawr4bebItZ:\\\\{swf30xz@aCyhb?af9Wz+70bWw*r,qWaUqeb7bas23Jxruqz/x698u26Wnms9*but;dm8bdl,eBaQxb6abau-|gbY/bu,eYaFnjtOaXsA9VuqmJ\\\\}?88bSazbE;ybIm0u>rZkNakuN9vbYa\\\\{u8uMrS\\\\{Z91|:pmbus-bwf;ppnH6?y7;Tas:?.cb/bQ7l\\\\}s/zb-xgbvtA9kuJ75b,vl\\\\}Ra2t>awbxbGa*4.9Yp>a,bybcy-b*b7b4b+\\\\{yzPavbEg2vZqA\\\\}7bGe71Wa18@,K:/p5nhbubQa=jcbXafw=aPpOa/72txbmb@\\\\{C\\\\{1bhb,bGa;,O9V0wox.Guv,IrEi/mYa>+*zLmo7<uBajbgb4*r:8bHtQ+4b\\\\{bkbwf2bvbl\\\\}*n,uznm.6bqnawRaDvCaubfbzn9qV4kbvbhb4eA2jbUn0*S5.bMjPmubq,8b"));
$write("%s",("|b\\\\}b8bi28b\\\\}b.b;p*bEafbFaa*+oxb6b/bQaQaS5,8Yn=\\\\{2b>vxn\\\\{bOajbvmtm+wAwYaQaGb?.2bEtM4KpmpjbfmdmbmkbO6,swbH,+seb0nrr1lFa-sDaYzvxp6I\\\\{/mG7vb\\\\}7tm0bfbfbibwb;5fb5\\\\{Xaw7fbhb6b4bDa3p7zF-04Q7Zk=ar7>qKx,8Pa9x-k**PaMwQamea2lbI2Hp/sFnbb+bDaEaU0\\\\}bwbababEa5\\\\{ab.p1o3bxbQ1tb@wDa8o5bkb*bwfusSfXr2whdns9bN-mzgxibxbwfebV-T-ibgbp3H6>x<x\\\\}gl7-mCa*w,wAr/btb>aF-H\\\\{K\\\\}xbzo|bn/,hxdWplpM\\\\{K2\\\\{o|b\\\\{u0bwd6/16h593yb4xWaXa;n?.mbVz5booDaPa4bBrM\\\\}|\\\\}.b=amtt.26EaA+ntO\\\\{csyb.bUqlb2b5g?njbR4vb0.s+Ua>ambR+ab1oQ6n/D20ofbEnRa2bv00o?amz/bjbFmI415e5?|zbF2\\\\{b<awbDa@aTavbbbgb.b,bW,5b;u23tb9\\\\}vb*bBa|bbbf2,3s2v*<wXak-bbFaZaY55nxbxbu4Va=-zbV*V*mb1oxbtb1o.ndbKy*,|,S5h\\\\}UrTx\\\\{bn|7pbbwvTs+bFajbTawf6b/59sNaTrzbibUe\\\\{dNa,vJqXp:3-w/bZ/dujbPnE-c|dbhbcbk1hnvbZaabUaWzXa/m,bcbxb\\\\{b=a/"));
$write("%s",("b8uabFa?.@pPaQ4Esk+hb1bXaI\\\\{0bbbybG40u9-L.\\\\{bUaCeogFak|Y-bvUai*\\\\{b|b02ibOywfMolb+b\\\\}mbx.bkbbb8b>,7b3pvb|4xbDao/EaArGojwhbBa@aSvabjw7rbbRah/Np=a3bdtAaybZaSadtwfvb,z?a.vF,Pad/Ua.vhb-bOaWzb+Uvxb..|uvpy*3bIxXaBvE1JssrGaL3sreuQ+Im=a.jl2jbOacb1bUadbIxiq|b<a?aDoybY/EgkbQoaoFslbYakmwbgdHqdbPaNt5bXaFaOaWawbFa4bWm=\\\\},|s0/bWu;\\\\}lbbbYaX\\\\{ju:\\\\}c0peXaBaVuC*NaOae3Ta<v?.0\\\\{A/ey3*5bXpfblr|b?aZs,b>v7x0bwfKqIq/bV-QaXa4bybVaNrW\\\\}\\\\{bFaKnebXa+d2b/|\\\\}b0b9bum8,AzByaqT.XambPu0u9bVa\\\\}br.cbEaGm:wAaqnAa,z|/H1fbmbPa\\\\}xcbbnM04bCacdBa5b\\\\}\\\\}/\\\\}l-lbwbPy1bZ/Bw1b>ox0v0*x-b\\\\}b@atbW\\\\}fdwb>aRaWakbQampTxWaCaA|fbPa/bwb7u0b*bebUv|wH\\\\{fbH\\\\{*bZodb\\\\}+8bFalb4bNaBa*b1pqv\\\\}gbqjbYa7z\\\\}b+bIu5bEa7wbb1nZaIglbGakx\\\\{bXaUtOa<a7bNahsZa|bWalp8uVahbO/s,5b*wG-L\\\\{J\\\\{8b.w,bSa?.V-@a1bl\\\\{"));
$write("%s",("1bvmqslbDw|b|tdbt,4pO//u\\\\{bmrYavb|,\\\\{t.b0b6b3\\\\{BaSa=aSwYaTaWwRaPhWaDzdbur+ucbmzft:tAajbdbRa3bep\\\\{b@|hb\\\\{t<a\\\\{\\\\{jq\\\\}yTaX\\\\{zrDaOp8n@m@al,6pXaZaQas-DoxbjqymFuQi2v\\\\}b>aqs;ujb*bzbHtRambWqUqEa7fQaYaWa.bSwlb1tAa8xeo*bM\\\\{Za5bbb3b/uQat*YaUanv1b?ax-lbtbhbjbybkuE.Kpn/dbUa5*XaPambgb++U.-b9bwqvbD.Ya@aVa7wwfWa\\\\}w>v?a3bXw<.;p=aabB\\\\{0m>awf>d=aFaAaSaWauzKnmb\\\\}bCa>v>a4a-,jtcy\\\\{b+,7bx.FalpMuTa4bK-ku;pfbBa6bMp\\\\}bDx=a<axbcbtb3pkb1nlb:q*bdbtb/e.t9nn|ib|,Ca\\\\{b-\\\\}Da3vV|=aQa9xupvzhbbb\\\\{pCrVazb3p6y\\\\{d,rNqMr*b=aYaRa4bdb8u-bAaXahbAa>aEacbXvZajbos1oNnQaYzOaRazbwbXqPaCeQr3\\\\}@\\\\}ybqumb*babSajbYoXaDaMv>aTa=t+bntIx;zZzorMr|b2b+bcbVw?|DotbLwzrsy6btbpncpNaybav2n@sOylb7whbFmAvMtcuZagb/bRa?awf,eiqEaPajb\\\\}*wbRawfcb7ttbtb2,Koxbyb3+as+b8t|bcjY\\\\}kbmbNadbcb4bio=aVaxbjbfb3bz"));
$write("%s",("bgb8bXazbmb,b\\\\{byeBnms1bjbbp7wcbRaNa=a,pN+lbkbEaZn1+.b/+Eawb/sSa>vVlWaWaqymyQa6+4+hr3b8b3b>aq+/bTaUa=aEadqQaEaAaVa=a2b5o\\\\}+9tEarxTa@ajtlmmb@apyOavzBambqyPaWa@aSaEamb:wOa.b-y4bL\\\\{*\\\\}Aaub>a\\\\}bSaBaFafbCjabcbhbab4\\\\}xp+bmbabqgUambSson\\\\}nv\\\\}tbw*AaquV\\\\{4\\\\}Ba2bYaAaib4uSa9oYaIs=aWa4\\\\}gxzb3babTrd\\\\}Ya\\\\{t+yL\\\\}bburgb+bYatbGpwbgbubEabbwbI\\\\{Rn:z/b-nYpSaDaD|Kmkbjtdb3b9bmb/r7bAakliyebib.bxdP|N|L|J|tbh\\\\}bbXa?a8bAaez5|=\\\\}ebcqPakbKqtblb\\\\}bmb3bku9tvbdbBaq|Zaau|bRa0b\\\\}\\\\}VaXaUaebIuwtcbBaRaEaq\\\\}-bexgdSa9wzoctSsWgzwluOq>v3bmbdbabTawbEv/bAaAavb:rQp,einfp@aaq<aB|@|>|judb<amb|dibValuOa2b?rXa>a.bWuab0bcbgbwblb*bFa*bQx=ahbxbstDrQakbguhbzrXaQazuep1z:vhblbep|bmb:vVa1bFaybfb2bEaFaeu,bRaJpZa1bOaAacbtu2bCaUaIbYacbibEa1b/rEaCaVa\\\\}w3bwsmb6bZaEatbwfjw@a4bCnwbkbPalbnp<azd"));
$write("%s",("jymq8v6vQasr9wybpxQaZaVaCaCnAa,bDatbFa=w/b|bubUaEaebVaimoy*bbb/bUaFa=tUaDartFaxb\\\\}g=adbXalbDa.q2b3nDamb2b7bzyxbPa-eTaOa0b-zBzNaPa>zjb<zQa9zDa5b,z@qzbNaEa|bAy<awfBawf0bZakbxuvbCafm+b,bHr2b9bFa0bDa*pXszbfbCa3bVaTaTaSa/bDneb/s3qmbubNsDaYqAa\\\\}xgbynVaupXaFySagsCyAy?y.bZuXuCaQaxx,bAabu1u5pkbnr5b6bctgbcqLm3bTaZalbAa>vvb+b5bebRaDa+bfb+qIw.bYotrzbCaTafb=axbabeb|tQobbPprtys,n3bkbcbSlWa=aSa.bRacb4agl7vAa*p/tkbFw8bDxMwEaCrmp6b1t/t*b/bXaab.brvcbrpXgWa7bDaQa8b6!![2aba!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"g3b[2lpa\\\\})1(f\\\\{#(tnirP;)23&=,bjbkb-fGa1wax/rabRaab\\\\{bnv+bib8btbPazbJwHwYvvx3b=wrr?s7b>aUaUaibzp\\\\}blbCq+b6b,babWaivNaef3mWm4w\\\\}bvb?adb.bSaCabbP"));
$write("%s",("a0b?awdSwPa-b3bMrmwub=u7b.bFaYlvbPa4tCafbiwgwPaTaCacbTaPaCavpdb|bkbpq0btbmeDawdlwwf-fwfVrlvab*bmbCaeb8bEaQaKnWaBabbIcXafbyb|tFm0b>acb\\\\{bib1bQa6b2b-bQa,b5bDaNa|b@akbkbOa-b6bdbFacbubmbXl.bzp/bBafbbmUajbBrcbDaXpubtbibWalbgbWabblbPa4anqQswb<a+ohbkb0bRaOaybUokbbsZr-e=a3rwfwb6ocbUaZkSlwb?aXaOa3bCa0bUaIcTf,bLf\\\\}b/blbub-s2bBaubWa9g8bibcbbb6bBa,bPaubybwfArub<a@aNsvbXa-kgbjb;s7bntqsgb7b3b,bfb8b+bBadu2b1bTacbFaEazb1bdbEa*b4b@a0b+b@a9bybcbOabbab5n,bbbZamb=abq8bwb.bwq3bYagb|b\\\\{bubgbtbSa7bcbNars|b7bUrubXs;pGfTajbbbEaJo+bXa3bFa-bwmdbsslm4r\\\\}bts<a.jri.bVajb>atqEiOaFambSaYa,bYaCaBaebRibbbbNa\\\\{b6bNa8b?a1bqt1b,bXsubYrXatbzbZcubTa4oibwfoiXaTaZqWa-b8b=aCa7b/babtbvnlqub1b9bUm8bIceb\\\\}bib\\\\}nzb>a;ruo\\\\}nznqrVamb;n*bPa\\\\{b\\\\{b.bYaVawf8b7btbzrKqEa\\\\{b8bvbub\\\\{b5bYafbEawfdn-b"));
$write("%s",("8qabvb2babybQa|bCadb*bAa-e@p1b|b8bVrMoWaqnjb7bXajbebPaXabb.b*nxbVaubBacbZa?aXgNa/bZaubzbeb1bcbjb8habibhbYabb\\\\{bwbyb=aXa\\\\{pSaOaBazbab\\\\}bebNaebvbTaQqOqtbmbqm+\"\"),\"& VbLf &\"(\"\"pebvpgb\\\\{bAatbdbub7bfitbTa+p5b2b,bQaxbNaVaDq/bvbvbmb+bybdbYaWgPq\\\\{ocb\\\\}bOalbwf\\\\{bWa0bWiOayn2oFm?a\\\\{bhp4bAadbgb,b6ban4bmbBa8bpivb\\\\{byb@aQm\\\\}bzbTaFa7bSakb8o7b3n\\\\}bVaqm5bwbCawfibFpyoZacjajilvnWaubwfUa\\\\}bdb/bSa1btbeb\\\\{pVa5blbxbJk2n8oSaFaebWaQa1bfbOa8blm.bOaib3b6e/bPaibUawbJkXaCngb0b|cOa4bfbabwbmb1m\\\\{b7bTaxb/bVakbNaog0bkbzb@a-bfb|b6bTadlib*b@a\\\\{b4bubabZazbUaxb-f>aeblbTaYadl\\\\{bYa0o.b?aebUaZafbQalb7bybkbZa4bZa7b-b=a5bFaPavmkb|ozoxo.b\\\\}bDa6b-bFa>a+bjbUaWa1bWajb9bNazbRaUaNa7b5gOaub3b7bVa0b,bOacoao>aNaAa2b@aFa+bWa>aFaAn+b8b@a\\\\}bTmbb4bjb.bqm0bPa,bwbwbGaVglblm>aib3mmbwmLm\\\\{mdbmb"));
$write("%s",("Vacbkb2bTa=ajb/mOaDazb=a>aubgnXaEaDaFa3bjbwfzbDaDa3bAa0bdbDa|bAaFaSa4atnhljl9btbbb|bhbDajbSa?a,bZahb*b3bEadbibTaab6bFa1bebnekbdb;dMjwb*bYa+b|bVaFagb5b9bTaQahb<aubJgWl5bgfPa5bzbkbjbibvbVaBa\\\\}b,bebCawbvb@a7b\\\\{bhbWe.bjbhbTa\\\\{blbhb>axbzbEahd7bdbCaEaybCeQa4bSa>aDa*bibBadb9b*b-bEa7b6bAaEaOj>l@aDkrk@lGlMjskuldkej8a4l9lXj<l\\\\{l6l;a8a.l3lYj2eVj7lVkyl|lQk-l<kolUkhkCatg0kWknlwbncOj2k<jplAkGkEa@aVj7klj/kNjLjTjPkNkFj4abjfl9acjdgZi/b-b4b/fKgubkfkj5kOk3k9kAa/fBkGeob@kmj9aEaOafj\\\\}k:kpj-a4iyk6k4kokfe:a-bfjSjvk=a0jKjqkPa/h|kqjojxkakck@a<a-bkjpk?jnkskUj-jIjik1j-aSgek5j\\\\}iRjgk:aCafj9jZj>aAaVj;jOj2cvjyj+jAa?aIegg/jJj@jHjzbrj,j>jBa/f.j:j4j8j*b=d,gpe5bxb5j4i3j*j@atg|jkjtjxjOa8azjSgsj2cAatgnj\\\\{b\\\\{jjjrjFaojmjfjuj?fij9akjHaggXi8aCa@a/f1bne8aej9f8arb8a8a2b4a4a3acg4aagJf3bHb6"));
$write("%s",("btgIhzbxbub9fKhWfUfSfmfqd/fld1bzb.b+ikh5iiiThAa=a?a3a8bLfAeSb3ihgyhzi-h?a=acguifhffYhTgvhxhSgkith>aBabggg?c|bvbmg.b3bJaEf\\\\{hXh0h1hihBa?arhzbIbKgrbehDfPglhSgjhDa2eghdc3bVf:bgg>g?f=fIb+d/ffe-b3aAaCa3aKa\\\\{b;aadwbdfIa3b1bEg,b|b0aAeob.hwhObuhNgCagh.f,fAeIdCf4dRgGeSbmhdgMgmfybehAe4digQgggOgBacgagvg;f1a4d1aOb8cubwbwf,bafPaofAfYe?feg@a3a1bdfwb+btg<fRc/b8befHc;a:b?fbeYeag|f,dZatg+gRc5btg/gMf3bKf|dzdVf/fwb-f3bmd;a<bYe:bYe3b-a?fQfzd,bxb2b2btb;aAeHdfg@fBf>f3a>a3a5a?fUcYe/fTf/b3b4b.b9f8byb2bZctb2b/fxb5b+b.b2b?aPezfIdxfPayfsfmfJbeeHaYe7fyeGavfxb-b\\\\{d4a-aYe.b\\\\{bXcMajaYe-bYeGeMdrfGa+bpeafYeGa5aGeHd6cYeyd2bzb;azb-bHb3b2bzc?a@eHeFeRaYaOaVafbVaibAeMd?e=e-a?a;a>a-aPaBaNdVaNaUa?a?aNd-aebcbTdvbpbEaOc7b@a@aDa?a>anbpeub.b+bzb>bMa0dVd<bFaFa9a>a:b;aZb8d+b+btb\\\\{bvb3b+d>b-aLcZb"));
$write("%s",("KbIbGb;aTd6akcOdNdUdRdZb/aMdCbKd6a/aIdMdId9cFdCbHd4d3d9a2b5a>d<d:d8dxbvbtb+b/bxb1b5a1a/a4dSbZbVb/a6c:aIaIbtb,b:avb|b+bub4bcb-badYcWcHaebdbJaGaxb,btb-b8a1bxbwbtbxbUa-b.b|b3bvbxbfbZbnb5aIb.bpcIb-avbocmc6awb-bxb6apb3c7bGa7bnb9cjc*b*b9chc/aObRbCbNbLb>a8a?a2a6a\\\\}bKaKa6avb5aJbVa?b7bHa=aGa>a:aGaCaJa\\\\}b-a1b.bybUbZb|bZb7aEaqbZb2bsbsb/aSbMb5anbHa6aCbObsb*bCbobBbNaHa3b-b|b1b/bJaNa/aob5a/a5aJa2bg[~ia3(f\\\\{#,43.3\\\\}ia9541(f\\\\{#X3~ma(f\\\\{#(tnirP;)23\\\\}ja7362(f\\\\{# [4Lma5904(f\\\\{#q\\\\})6j3bh4Tg5Mda132g7Tja5683(f\\\\{#&[2iha=s,y=z,s6[\\\\{8Qea0603+:Vba0-;\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'i6[Y3+|8jk5[-;Hba76?Uca560<a7>[u8[6=iyay,]99999[gnirtS wen=][c n3aea\\\\{)v]y3b&a(niam diov citats cilbup\\\\{RQ ssalc[4Lba7@DVea9493$?[h9Uba3~@Wba3~@bj:[9a& cdln&&&&;maertStnirP/oi/avajL tuo/metsyS/gnal/avaja:"));
$write("%s",("b&ategn&&&&2 kcats timil.n&&&&]; V);=:a;3ecaL[I:aD:hha dohtem;3a/4nga repus~3acaRQ83cgassalc.|>[\\\\{:Rba5>E(\\\\}9-ca14#:(i6[\\\\{:.oa(=:s;0=:c=:i;)o9ajaerudecorp>=Mba0$Ma>=Qba9-R[PF[g5Qca75.RUza1251(f\\\\{#&(tnirp.biL.oken\\\\{,9bianoitcnuf/G[96[A8[.3cba1BNWK;[qa(rtStup=niam\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'tni[>Nx8dkawohsn\\\\})840h;\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'MJ+ba8~7Uda332Z4Qea1918c@Xha=q\\\\})486h6Uca148GQba7f9bta(amirpmi oicDAx\\\\})42QIaca3Cl3fpani;RQ omtirogla?9Ml4bk6aea.tmf>Acfacnuf;t4Tdatmf[3Ugaropmi;|Jafagakcay>Mda115)6dbapu6Mc4bba-X3Sjatnirp tesu=MyIaca(n)BQca725:a#a,s(llAetirW;)(resUtxeTtuptuO=:$5Mca36)6ea4RdaS CZ3M.3aca&(X4Rba [5[[5SiaRQ margof5O.3ajaS D : ; Rm5Tba\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'X3Sqa. EPYT B C : ; Aj5Tka)*,*(ETIRWt5UhaA B : ;e4Sba [2cj5Vba:a4(+3[+3wda(nfKC&;Ya|a(etirwf:oin\\\\})8(f\\"));
$write("%s",("\\{#>-)_(niamp3cpD~ka(f\\\\{# cnirpP@~T4ahastup.OIVO,FLataM diov\\\\{noitacilppA:$[cea[06xE3k75a*Mcpadiov;oidts.dts 5Ka14\\\\{kaenil-etirw45lva(,\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'s%\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'(gol.elosnoc;)\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'K3s[2cya\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\' nioj.)1+n(yarrA>-)n(=ff4kia!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\}54,1\\\\{.n3cja# qes-er(YRdba&l5rba!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"$Sk$3lo3r33tla1% ecalper.S4l(3cs=gsarts(# pam(]YALPSIDq6cua!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\".NOISIVID ERUDECORPU3kma.RQ .DI-MARG~3oE3dnaNOITACIFITNEDG9dsa[tac-yzal(s[qesod(n6apa!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\");\\\\}\\\\}!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\");\\\\}/****/e3a\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"),s[99999],*q=s;int main()\\\\{int n,m;for(;*p;)\\\\{n=(*p-5)%92+(p[1]-5)%92*87;p+=2;if(n>3999)for(m=(*p++-5)%92+6;m--;q++)*q=q[4000-"));
$write("%s",("n];else for(;n--;)*q++=*p++;\\\\}puts(s);return 0;\\\\}\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\");gsub(/!/,\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\",s);for(print\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"define void f(n)\\\\{\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"00g,\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";for(m=1;m<256;m*=2)\\\\{\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"00g,4,:\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";if(n/m%2)\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"4+\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\",\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";\\\\};\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"4,:,\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\}\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"389**6+44*6+00p45*,\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";++j<=length(s);print\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"f(\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"n\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\");\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\")for(n=9;substr(s,j,1)!=sprintf("));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"%c\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\",++n););s=\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"4,:,\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";split(\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"145 160 17 17 17 23 252 141 0 46 125 231 229 231 250 151 243 243 243 231 231 207 159 63 4 231 249 255 191 225 17 127 206 103 5"));
$write("%s",("1 57 152 37 255 57 204 230 103 48 79 159 159 151 252 231 51 51 57 193 47 249 204 230 102 115 4 251 190 249 243 207 57 206 115 158 9 231 57 156 206 102 9 193 48 96 22 236\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\",a);for(i in a)\\\\{s=s 0;for(c=a[i]+0;c;c--)s=s\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"1+\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";s=s\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\",\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";\\\\}print s\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"@\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\nquit\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\}\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\")');\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";FORiTO UPBtDO INTn:=ABSt[i];print(REPR(50+n%64)+c+REPR(50+n%8MOD8)+c+REPR(50+nMOD8)+b+\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"J\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"+a)OD\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\"\");end;\\\"\")\\nsys.exit 0}\"\")]]></xsl:template></xsl:stylesheet>\":s=\"   \":For i=0To 7:s &=Chr(32-(Asc(c)>>7-i And 1)*23):Next:System.Console.Write(s &n &Chr(9)&n &\"  \"):Next:System.Co"));
$write("%s",("nsole.Write(n &n &n):End Sub:End Module"));
end endmodule