module QR;initial begin $write("%s",("Module QR:Sub Main():Dim s,n,i,c As Object:n=Chr(10):For Each c in\"<?xml version='1.0'?><?xml-stylesheet type='text/xsl'href='QR.xslt'?><xsl:stylesheet version='1.0' xmlns:xsl='http://www.w3.org/1999/XSL/Transform'><xsl:output method='text'/><xsl:template match='/'><![CDATA[write,format=\"\"%s%s%s\"\",\"& VbLf &\"(\"\"\\\\write{-}{txt}{(\\\"\"with Ada.Text_Io;procedure qr is begin Ada.Text_Io.Put_Line(\\\\\\\\\\\"\"print\\\\\\\\\\\"\"\\\\\\\\\\\"\"STRINGz:=REPR226+REPR153,a:=z+REPR166,b:=a+\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"2\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"+z+REPR160,c:=b+\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"8\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"+z+REPR165,t:=\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"write('implement main0()=print(\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"BEGIN\\\\{s=(\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"#include<stdio.h>\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\nchar*p=(\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"Ra#include<iostream>!nint main()\\\\{std::cout<<(!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"class Program\\\\{public static void M83apbSystem.Console.Write(!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"let f(c :Int):Latin1=if c=127then!!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"!!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"else(string_of c@!!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\" g caffeine !!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"@$3kEa!!!!n!!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\")@f(c+1)in print(!!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"Quine Relay Coffee.!!!!n!!!!nIngredientsq3aha!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"@f 10U3cgaMethodz3c#a);let g(String ->[])!!!!n[c;t]->w4edaPutY4spa(int_of_char c)05auainto the mixing bowl|4ejag t!!!!n|_ k4gtaLiquify contents ofE3oeaPour\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'3w\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'4elabaking dishv6biaServes 164doain g(!!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\")))s!![2aca!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\" [2bo3cparts(nltnirp(])]v3cja.NUR POTSp3cx3dp3jba!!M3dp3df4fda[))j3ci3e,3cp3l[2kga\\\\};)06xu3n<3|ka)1(f\\\\{#qp]\\\\}13$fa3(f\\\\{#+3~ba7+3&ha51(f\\\\{#.U3\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'M4&ga(tnirP%5#ca72U4&ca36,4&+3,h9l,3tkaD ; EYB RC73(da,43.3\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'daDNEZ3Sda. Ab5VeaPOTSc5Wb5TmaRQ margorp d&Baj4ObaSj5UV3Lda721W3Wba&R5MY3bgaS POOLl;Vea\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'&,)l;Uga. TNUOf5Tfa(rahcp7Nh5cgaB OD 0o;Uca&,u9Sca)Av:Wq:UiaEUNITNOCdMaca01t8Um8Vo7O~BceaRC .b4Ska,1=I 01 OD9FWcaPUc4Ty;Sva;TIUQ;)s(maertSesolC;jSms4<la552(f\\\\{#n\\\\})6i3ag4Mda115X3Qi"));
$write("%s",("a3201(f\\\\{#KT%z7*ka402(f\\\\{#mifb4Nea5904\\\\{9Q[4bba+[5U%a315133A71/129@31916G21661421553/\\\\}4Tfa(t+s+b4T|8Tsa(amirpmi oicDAx\\\\})8;6cgaCx\\\\})69f?\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'DZ-xa5531(f\\\\{#ni;RQ omtirogla87V~anirP.F;\\\\})1+69%%))n(tni-i+512(TJN\\\\}4bbaw|5VhaaepeR.SZ9UbaWY3Tea=+s\\\\{&>U#AU$ENia918(f\\\\{#\\\\}\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'DOea91339=Tda760:=adadne-FOea0471f5T|a36351(f\\\\{#PUEVIGESAELPn\\\\})631w3a[@Qca36\\\\}5aja1,TUODAER\\\\}4a58Mba5\\\\{Nbp5Pda110C?b\\\\}aetirw;\\\\};u=:c;))652%%)u-c((||V;Mba7#Mb~5Pma99422(f\\\\{##-<[=Nca97c5Ula7742(f\\\\{#||ij7Nea5965=;Uda707i7ahaBUS1,ODh5Mba7mAVea59395;gma)3/4%%i(\\\\})882:Vea3060~5Uba3d5bVWOba4\\\\}6a2EQba4&8abBSca111:abBQba56<aaBcNa2=:/t;2%%t+2*u=:u\\\\{od7 ot0 yreve;i-=:u;1=:+i\\\\{od))1(evom(dro=:t elihw?s;)s*0>Nda9914?aW5Qda758:Bb/>Pea7881g5Uba3s>c0>ci5Mda"));
$write("%s",("659z?Wba2(Ybfa\\\\})293PMVca97PMbqadohtem dne.n\\\\})82OMWca34OMbmanrutern\\\\})409SLVda768D7aHaV);gnirtS/gnal/avajL(nltnirp/maertStnirP/oi/avaj lautrivekovnin\\\\})23*LXca35*LatHN\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'LVSFZea6962.Yacb\\\\}\\\\};0=q;)]q[c=z(tnirp.tuo.metsyS;)0(tArahc.y+z=]++n[c;y:]q[c?n<q=y\\\\{)0>2%%++i(fi;48%%)31-)i:3c&as(+87*q=q\\\\{);63951<i;(rof;n)rahc(+RNN$CV47Zb4[b4[kBVca16@=Qca33l9[b4[b4[KBRva941(f\\\\{#=]n[c);621<n++6>aqa0=q,0=n,0=i tni;XLNba2%HW/7[b4[uJU(b8932(f\\\\{#6aeeicpbocJhLfbR6g3b+bwb-e62JaMa\\\\}bJaLz-e-bJaJa7zJaJaTaJa8bGn;a8bt*Ka7W@BH+l0Z?8pbR9bKa7WCPTa7W7W@BbR@AJaLaJa7W8bbRd4cqa8bbR4bbR:b+b3b+b&4cgal0JaHa#3aca@Ak3aGbJaQaY/;a7WUa:aUa:aGnocXbddxepgXcVcScQc/aDg|bb>IcncDcZi@c|bKa<c=a0c@aEa2a;c9c7c6c4cAaGa?aJBJa|bxekcpbzc-bCdlepbocHazcHapb6a6aIc7e=a-awjed3bHd6a6a=a-a"));
$write("%s",("?aY.9i3fdb:e7apb.6FeDeBe@e9apbGeEeCeAejd1bMwYb|dCboi:k7a.6,h*hMawjedvfvbJa>a2a,g*g\\\\{hMa?aY.CfXbybvd6a13i6bHdtby0vdie=aSeRaX<bfX<kb;xttSe?hqe7b5aIgjcYcWc6aSdwdegSBBhMbUfUfIb/bHdlfjfug-b1bK3Hd6aSd?b0d@jyb9asi6aUj2a5aqifeefdcMh4ajcJg|b|1jc?a>f>hz6ak3aeari<bv6albkf7hNdniP@OrBb@bB4;adghf?BpbP8NK>b7;PfNCyg-avfvb?a>f2hCd0h:gEaAeyhwhAaSf9a7btd-a5b@=whAa3a=a9a7b7ks3g53eea3aAa73kI3a53iha,b9a7bn)3hxaL0Jh9a7b\\\\{L-a5b.bWklhvg6[3bk3agaKiLE<eq3agasbwhEakA~5>/fa(f\\\\{#ac7an6auaLgwhCaRf6a?h>gOgKh:gk3ckaUhuh<b3c-ar8cA7cda/h?73aK3d-a<h:h6a<bxfig2oKb2a=lSgPh8fwbXcjc@aCcVc6a,>a&aub5c5aye=anbSgybph5a\\\\{e6a7bJgHawbXl<bsa-b9a9b9adhSg-a6a>ao3aea@a@aq3a)a@a0c|b9a0b9a@a>a7a6a@a>aIa|b>d9bJa0b-3a#a-b9adh9a1-Ja9bSgnbJa6a|b5a,bHaH4aga,hJH-aN<a%aVt/fVt/f6a8b5a1btb*e-a/w@Z.bbb-a\\\\{3aba7\\"));
$write("%s",("\\{3nka=ljdEfNHHd~4aua8b9a7b5aMaJaybfjWQ1ca?awaHajgJa,b5f1cJa-b-a\\\\}c\\\\{cs5a)a<a2b.e|bMd:aJhJaub5a-eMd?a,bSBJa3bjc[7cgaIh3a3b0<e;7a5eThRh;aYcWc=l9*,eIi9i1jmkyihjWj*cyjrkakl9<kBh|q+z1bqA77gbs,0bxfhxWkjbSa,b<olhLz\\\\{PMns\\\\}DN@/B*uIbbkbJ:++DLEalbV6++zbYaKu2bhtjoI?|z,bqA-l.zJd0t=a>a;|>ax59x7y8mCqdbJd,-bb<<DaQo;<fbE>>axlxo9*-lYaEmJSOrKnVxc:@aLA/m-qgbebj\\\\{/5=a9sBx3Pb:.J7y0bu>VXO29t.bO?.qhbTa;>Bas>\\\\}<7.\\\\{wqyAaNq5bVFfn@>7WJH\\\\}qZXQwjlJsKnBx--lb5p|9?a4|mbr0zEw4EajBi<Oa?s@yTa.IExq2mbCl,bWa?|wb3y=3m:bR<aTaYvkur|0uss?oumUpw1eL<COaB:<kJpCDGl\\\\}?/bHLLya115(f\\\\{#(ntnirpn\\\\})652(f\\\\{#<[$n4/TdYWIu5b+6/uUr.nO?D<Rp*1Yqz-xbnlxZnnQ\\\\{9spdKU>xBa2d@aeudKBaNrUrsOx.B/bnM,\\\\{b<a,bVoOmMvVaCaDq+h\\\\{veHyboE;r6qbbv\\\\{Hybb.b@:Ip/bT,MV0bzxu-H5klwqGZ<ax9H7jbZl|ztq+bI+wMibYkQ\\\\{vbPme*Px"));
$write("%s",("onWICtd;nnebG7vxJSEay>>qqKAg+Mnr=a<aYarq0J4;7DUVS>uUHwVmfbfl|z,bxlLeh=Sa,bqAP>FaqKlmEadvmrT/:n*b\\\\}4*sb,=k;kh?5>/:ZLPxAkIhhb@|ubXnb,iKGl<S>aN>Ryn<r0a7lm@7xxDsupp;fqvm>aWa;w\\\\}3adbM?qB7>9*<e0uomSa\\\\{pjbZabPPazEDa7y1Ejb|FSaDa5/DavbRmQMM:ubmy>ee=3k5/YBHd-b++u++k-l.nV.+k-l-uc3aua.nvbIu-bL=++lbA@H=O=k3cPd@+G=t?D=kCA=k=TpylvEtsiAYBNl5nSakbSr|zlm/=Qxyk++<kQa.k,bkM\\\\{<Ea;FfypyUa=.6\\\\}++@=Qx/myv==NZ@Ua7,bPF\\\\{<U4MeDDSaKW@/DDSawC5bDaY2WVAa-u-lYa=;G<zxCH7bpoE,Da7l:?BaE,am.7fmZaQ/9*Ca.za4.zVX.zQx4<2<WVAa.n@|ubmnQDK/yo7b<?DatN9Gbv5?w<E+flWly7fbD6u,l.+kl<hb+n0u1l,3=aYa64a\\\\}k\\\\{5khbA6fmUlWD>adbgVE/ZxGndl4ldbytV*9;XlDa?aDadbE0CwZx>a3+@;hbTh0u<aF@wbSa|qhb)3cgeytxoslx5iK?++;Il@7hbK+q2=aGndlblhb,wt,NRDa3yn8x?E>L*x-DaJL\\\\{u?zym*eMulpXQX:2yV:GaA-8l=\\\\}xfabPl-nrsWz7buIjbvb\\\\}"));
$write("%s",("xIVHGnp>rV.nFhbNlDa?z=:1bP0hbx-A|nvS?dbhbmnupyb/bWL\\\\{9@a?+J>*b.bnIngNaRars>abb9ptb?wA9crmRW1>xAEThVx<a>aE\\\\{?a6wIlp5rs>aLpeb|q,bX7u,4QDaR*,kMu>\\\\{c7VrSaYaYavK,b@bS?nvE/abeb@k\\\\{b?sY1u9KSYa;9bqozuWebXaCavb\\\\}x|vJ<P-A|/bbguq0bdFebub/b=aq0mKgBz+rmgb.LWo<T@2fqU3?eaWa4OW3orfBom7ZII?KF\\\\}5om;n+bmbNwU;RydCbRN/e3Vv?vn?KOUK1\\\\{foAEvdhbTap8;>jB4nVvX>@=<rVvqmE\\\\{p..2/BcO8w@?jwku8Mo;kz*s\\\\}34tSGhbE/.=H1P1u5L*8cKEW40qUasmf8JI+@.Cu5wbwoJI8bNm2*-9V,3/X<6bxbYV0,Cxvd1bygkb64jbCl?akbe>-r@aS+tb3DlmW2IRBbt1tbAMc4IxnnLf12Tk|mx\\\\{p\\\\}M><orGgbEai*Yaj3vb9*mrFk2q8bh;:dubBb+qb>Ca|YOJF\\\\}3ns\\\\}QUi9PnYapG>a,b+h\\\\}DRa6bXc8bUr2/>?jwaoPzqHr\\\\{glUkCakqebAM?:mNZ\\\\{tV\\\\}bFDBa<tyb9bYbwXybAXr0zse3ybBa,e:\\\\{6rWv/BFDtq;tXa7zMs\\\\{OyNayMs\\\\{OP<U:5C?aoqGk0y8qLz\\\\{WH-U:ABJL@k>60>U:Zaih#3cQlPahui"));
$write("%s",("lDa*<a+ax.xaqmrr5p5Cq3yS7pm\\\\{biKdubuVCih4bmrWqWOWI-Liu9tCakbNCe?ozdv9*vbXBks9tab--;F1@TmCtxfab\\\\{<8bfCTaHX2dwuxfRv;xWahfxfRvUa0o/bYa4MSX2ASa=3z/kbEfArvz|KpNQDE6t9\\\\}b;@k-MwSGzbxM8YeE<vKqZXa,l|BXJpebWn\\\\}CGPOyU\\\\}M2@aAmnymbcbdHa,yo0bLohPb*Dtcbyb:mM7ctFakbxvU4+7NnK5.66nnqhb+q=zT,KzlrmbgUisVa?apsvOlbbbWaebM*QafOJv.P1xRyoE0bKr<rRaRaHxFz7b=wCDTzBa7bY\\\\}*+<DE=\\\\}bPm=3E>Ya+DGaIGz\\\\{9*qAJ-lNub97P8KuGnD.P8Kok=?u+=iYJ-?w|+<,OM5bg?G00\\\\}Z\\\\{c4RH0b6kv\\\\}><ihtlKKab=aT+j\\\\{>FhboB0Abu4<WsWapo/bNyLvXaK.8b85F0.:bpabphZekbHrGP:sNf=afO,YQp\\\\{bLxUa-+<xnHXoJOC5MmqBFhTaW<YnHyG-K.0bXo1sMZiHy|LxG=\\\\}DbrWZ3pXa@aR+cLao6L3*qByBJphbi5abcM\\\\{=wA>a4zVH5p606dGP*blb.b+F.*t*OyVa*jwJBxXEzQT+/wNX-wqJlqQYzux0z?NCkZxb2q\\\\{dG\\\\{KU7b/05w3n9bCb.m<8dukBImUaOth/mb>70b.toYJ>?<>,FaW?|=lbvd8b?s,YOr"));
$write("%s",("Vac+*b\\\\}YXx0p9w-bq0KnJLbMVxapCzvb=Ylb7;Ra4bK1wrIdRwG-xAkbAAP=\\\\{b7bJnQ,dptwn?LkEsm:zbtbx>+U.b0bys<O6ba@U;c4wrAaxfpA6XEaA@85p|<tPacbR+abCaew\\\\}+UH|s+bUavrt5M\\\\}\\\\}bDavL.mkwfs?L@y0umbzkVmM.CaZsZaZA10<QF.Vt:M.3T5ab>;rAtvubl+0Xy8q5Pa\\\\{bsW9.Qa\\\\}bfn;nyyLNRN?aNa+48\\\\}HrUIIkfbto@/GaaAym4qumc6F-;:0bjb4b*blIl+lzaln6xh14S~la(f\\\\{#(tnirP;hT#c1(f\\\\{#@<tTnxlhpis0Tb30pqyhltW0*<eAadbj6=0Nvgb+Bh+l9BAAg9b+bPa,w,bJC?L3+ag7bst=F-bTzy8Er>3n5fnkxnqZu,w-n2HSaOo@8gb>86bezczaz@>;Erq;2K?AjN:2HPam49uY4:=/b.bJnw1;VqUtQ-/w1,RT4>a*TY8OJ9*\\\\}PThPDRa0kUwzbrE+bxwwbbuebFDI?Z@ubWwWaooBAeHGad2<V:LIz,Uvzb2b3>tL/jzw1/b|4RyBN:w7m.btbAaCvs|zb?S8r6Lebj6Ua@?mb>?jb:KX:cq+UKtEoUaFa2FKdn?H1@Hk5;EopCz3/vz?aUnRP?<zb0bJCi.9bWa|bT,GwKU:?IuybxvTecgLoJxdb>nx1;14?T.@+tbrpisGoxf|bN3Yz4?CbSw,wx0ttC:IvWarE"));
$write("%s",("mbduDPHBTaMrQaxb5dbb6bZ7kbSti@4sW?gbYa?u6b>awb9*kbflC<C:6r9mdt0bQab>kn6bOaZ3.L>EQ\\\\{<o41Sa;ERkCy,?u,r|Wmtr*b9u+sJpv|?aSa@aS3W|Y3|K/\\\\}BfWaI-7beO8qKn3T,bQnvbt-MdWkEes>hb9b4bF\\\\}fbcb*Evl-F>IMvtoFkeH5.vb3t/B7k7kBq6dpNW6s9Bx/:WaEa--RaHrLxPlxfJSG-rrz+K.n;g>>BWaWpyI1uBG7tQa,bjbCHX=8rWlQafbnmc0Ftdq1bCawbDahngbmO@22A>q>EHf\\\\}bNIUaB-BF7*BE+zIspNSzDFKF9*hb5bkxun|p8bgD8b*E?aVQtq-nI+zvm.?0pyrnab3bQaB>+qP\\\\}P+P-fbcK|6m-nRs7SyHQhb5-?aTzVa-OCaPaf1:w*JZaPa--BNT>MoybCENfQ-*z0kvxUaM.mRun\\\\{pKo1E<*GCSyy//bOapscbQynHS3P\\\\}KQP-N-f?Wam.|pXo-OzbM.Wa1bAaHxUa;>mb0kOaFbPKU++b;6CaBN>aGaJBabG|R26-sp;r5CoMEakuNablD\\\\}VwiQZO42vGY\\\\};:R\\\\}WaYqMIkz8x1b/GRuVa6\\\\};F:0@\"\"),\"& VbLf &\"(\"\"ao;4bUnn2yb9*cb>I|savbbr|ErFa,.Dm?.Oa8Mmboy6AZ/;vTe8z>m/0,?<aVaOv@ahyJO*D3:Z/Raa\\\\{X\\\\{QDk0r@v5+lkz>ahb3b"));
$write("%s",(",lqA6sqH8b1bTpVaRa2bMwNa?aibubYa,t*t><HvXey7V/l2YnE|anRiZaUa-Ldbybcb>/HIo:Ta2\\\\}VaUaVx/mHdGHTnb04m,AGaDAID+bQIWavb=zSwhb?a7EJumbx?n,RaPOSanndKAa-Ohr?9.JgvWaWaHrpKOy>>Oawb/:n*SaTe@.v\\\\{4bC.yyB|MMq0Va6wR||Akbs4km2N>u9*9t3N4LD.Vm/LWa9bQa:w-\\\\{Sa4b>mRaOxG0jbYant.bvKE\\\\}4<N-H+FaKx942bn?ym6/Ra1bduKny4>1t|7sXs2biq4=vbn<<a+qp:*45bo>xfe,1bJCRFFa+wiqlbebcbssNki@kbe.>\\\\}h/ulDx6v-br,qAkmubW*L/bA6b3rKrN-Ta5b;6@txv*G7bd8xs1yt2EaYaH/:sXallPq/b1bX/jCTA,eSGhrHm@l/oEabqAqup*\\\\}j3eL7G\\\\}bxE|FTa|m+bSabbYa+bEa9r?\\\\}\\\\{=6rjxYvUlOqTacbzwji+?cs=lCI\\\\}|fbRafM=\\\\}yb@DI5mbt@FLy3ub9zAaon1skn=L|u7GNa8bumAwZBAAFka3Ta?ac6KqGa.Bd/H-Y:m-5b>a?Hhb-bfo@aI?;pbbxbmbZECatbkbZ<E7l0kn=<fv3bDx*y\\\\{baoL*kbYrmv?l\\\\}bUa6bJrrt-emJ;vmJE/Ua\\\\{q9bGu5eonzyOaPambgnGa@g,3C|xbJ|G-fGsqNaxfOaI+H:Tz*y,3Un5CjJw"));
$write("%s",("5Qafm\\\\{bdbIzXaU>>t@peH\\\\{|DakmnmRJ4b3/kG@ouIgb6d1bR=IuPI3bKF\\\\}<bu2ASzhbBa@a?wRa?F9*gr?|OJ?aRaxbAjhrQ,W?hpgHMsMmDp|uwK.r5Jm3Uafb?|Ve3bebVa=axb0>d7=.Sa=a+bXo8b5JRilbNa\\\\{:g+b\\\\}.bSa3b\\\\{b-mIJ0qvk0kb\\\\}XeMJwbAaVliz/bBJs.Kvft@oSaFJpo?w|sz3V6K<y,p|OaKnYzH0o:0k@a+b8r>kg+.7+..7yw.cn*jbl\\\\}<sPaOrbbkF1<er7l4/bb-bWzy5<aOa1bJH8uHyNaBbts2b\\\\{ko58r7yfl5sP+>b6w4bBwNaHr;qFaJ./brlfbjbDF4p=a12mbWak|hbAai*/w3oVtL,B9BpYHybebBa.5-slBT/HA;6|nKnS7Za3|wb0*2b@aPaRworknj27mwHwb3bClCqCa>;N\\\\{xbertqtlHuBg>aLzkp-m?aVacuns=mTz6/*b/|ZBewZa;n/\\\\{t-SmBailTw,b/bl.Ra8ktb:-bv3b2q>7/\\\\{DaNab>/bybWa2bjC5/x5+b\\\\{HHD:m1/W4X48b0*7G5bSGVutool\\\\{HVas\\\\}kbY|7mkb\\\\{vBaVaXoVo:5Aaq;o93bu*hf1:bg4bBaYakxZaH5ab0rapmbb>@tTa20W=7A\\\\}b3;Y4VEwESaK3bt>;xfxf9*<uMfupwvk.7+cvFoB4t6*C=a6oYa/ov1FaRFupuqS+f1x1\\\\"));
$write("%s",("}7jzKdSk;FMolbWalm\\\\{|ex:o=4WabbrGzb5CQaDF2bjAtb1@/kJ:av4br=3;Ya?<Xclb?zDsT3,CPmKoWw4nZlVa5bPt4b\\\\}s/p3y.nmbtqX/Xu*wu.VotbebGaO@Cacb9bPatblbEa>a:z.mW|apu82bAa;n=nu;|p?aGaYCEaUlAaL+ab34iFD.Aaq\\\\{Ch1\\\\{fbmy9s0bwbc<<9ubeFcFTqwyC5TEeb76h-pp*A\\\\{mkbwyCaGu-oi@XtTa9*f?Hu2n.bxbZ\\\\{0tkiR8ftt/vxZaDa.b.2eb3bvs5bVawbR2i*?:y<Pmx-0slpxfzbCa\\\\}ns?@amb6b?+aqjolbO7Fabbubzvrm|+2bkpi<=a7A*bbbXa=.6mW?HyUn\\\\}bjoI.QaGa4vasr|<aK-Ko\\\\}b@o;vNa*bu9+lbtc/dhE\\\\{yb,blBVa\\\\{3wbEayz*eI?JdVvZ\\\\{Qaxf+=/BauUa/k=an5Iy*pW6iuPmfv.:fBjbAatbY;Iv/k1b6tj\\\\{W.lDzviD|uQuZ\\\\{>aW.2b\\\\}bgbh=upMm2b12r\\\\{<tv18bo6oo2bs4Rak+tt|0;z9*OaY.Bg|bI?,3;z+b*bn7Vaki:n:d78Ba>tVans8/6C\\\\{b@a9mQkRlFxbz,b.bN/n,*ng4NcY|P+cq4b>a|b7<S,inybTa6bA,l>s\\\\}Tngbis41Nu\\\\{7FaXm,b@ae?+6m>YaAa|b\\\\{0;z76BaEa8bSzOa4b1y-b,l@,SuTA<kk-y"));
$write("%s",("b|A=ahuxfTml8W?lm-:bzTa8bfbFagb5pL*r:Z2rma|7bo9s,;n6bEa?axfwb@ac+\\\\{bZa*<t?xfn,vba4\\\\}b-x\\\\{bCl..1\\\\{Pan9wmI.Apwb\\\\{q-bFk=w*bdbA|9lgb-bjtybbb2br0*-w4|bZ4foiy9*>mHyGp2bjsj66wZ\\\\{D/9p;rUa*bzbwb\\\\}bXh4/@sQnj6o><a-bXaVnxbZ2N-BaJ.;r1bbbOxmbG-R+Bnxf6r/:ybRa7bubaqouY\\\\{P+ub=aw.52XajAW@\\\\}bNaM@*p\\\\{@3l.6aoxf\\\\{bhb*@rmLss|b*ib5pRw11xf5b?<G7xbcbrn=@m4jbeb:y1@|14pEa,vrn6bu>W2WaOn8bClW2+=|nubzo9ykb5ku9GpvrudjbBaV3Oa/bP=Bu\\\\{ppd7bM;|bj@ybClhwanw32uPakbeb4bCa:?js|gp56b.bE7Oax2Tq7b|+Tp|m9b1b9*WaYa,b*bTa+/G7Qa+e@3Yk4?Emn3BhVr!![2aba!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"g3b[2lpa\\\\})3(f\\\\{#(tnirP;)23&Z04bs95b|zNahl.bwnsopxalBagbXo8m7.x\\\\{*70o<v3bYr5bib4/Sa"));
$write("%s",("Fa8/dbFarqlb6bZaZr-/\\\\}9GaPs.br0X<<a:k09yb4blbm.3b.b|gct.7Xarly4A,ibabdbb/bb;>F\\\\}VawvlbTatpv5t6>aYaIpJ=ubrpjbVaAaD\\\\}vxSadu1\\\\{Vvb=<eDaw4Vb|6mtlbtmN-*mOk@aZp*lWzp+OaFaUa,bnumbOvPaTs-95/Xa,9.b8bl+NaXa46>aX=Easdn<2bY1fbJ<YaAwIu8cp5J=kb@+Ox-b9*Va,b<=Xo46um4b?<Uaduzbtsip,bCt.bp5OaSs0bJ2>tlrRam;Aalm@<n=WanvebMn-bZa?a*bkbfbOaSuk,/qHzd=+0Ls9b:o?u8v<a9b@/xf?\\\\}rt|blzrnvb-9=8Ua2ulbw8Oa|bSzR*U6?a,xlb\\\\}bUrl6N4fb=akb-uNtfbfb,lebOa.kcbOa8bwb2bibAak5p79vfbebPxRamb8m2bio?:+bUqs|kbLo<aSajb1m1gyzt6yx8uy,BqHf64K1jb*b7b|k3r|k8bAjkiFsDsh-tbWncwR;<e.zBrd-.bSoBt?sCa<a\\\\{bF;4bK-9*Su@+M.BpdbFm|b6qw80+nr?**bNa=nbqwvXa2b,b2be-2beb\\\\}p-bTakzZ\\\\{n7Fx43Z\\\\{@7@jkz8bek/v5be-8bWbOaZ\\\\{kbwbWaFa.bUyq52qinMmX:46ps3bS+\\\\{,E:;nfb5bc2C\\\\}Qac/@yps*smmpskb>a.bcvkbdbcbj/rt?zXa4bvb,3jb\\\\}bcs57p"));
$write("%s",("3RaRvx/:dg1Zl4mc:kbjmRajbUa|bAabwBajbx:kumb*p9szbR\\\\}?z3-T.6bvb@\\\\{Aa0b=ykb\\\\}3\\\\}bwbF|Iq@a+q|,IkcbWa3s|rBq:\\\\{ylwl*bSa\\\\{uulslqllhJdgb6b2ukp9*u,+n7bT5gbl+=aTat.@a0p>skbkboqUsF8By|bZwI6<axb9k7k5kYakbyb50NfDad5=agv1uxbPtC\\\\{Yamb0bvbz+Hf>as4jlvb5\\\\{\\\\}rjb275t3tppi0HyM7ewi*B4\\\\}bJ8ub|qlrGl\\\\}b<r|bAwt/@a6bWn-bF..bNaoz*q3b\\\\}x8bhbH1b\\\\{tdhbKm40C\\\\}>yNaTaByJi.7P16btbO0Z|2y9\\\\}\\\\}rAk++hu45>,dbxbE/lbD29bcbprubg1ibxbxfD5lbi.5z3zs376jbb|f,F|Rc\\\\{bWwZ\\\\{Cahqdy9b-bAaF|G1Ms8bK\\\\}vbOp9*UaUnOaYa\\\\{qPah/0b+bwpOaPn5bn6|bFaF6PaFxXa?+=a*rH6Tazb/kiqdbb0Ra.b=aXatb4b,u\\\\}bEaointod1b@a.bk5EaVvgbAa+bNy4jR\\\\}nnJ2|b-mTa=a\\\\{bSaG-w-Eh.bUabbPan,\\\\}bjb54ubHz;mEa*b4bPa>a?zyb0bCa|b?oZ*>k;*vb,u@vbb+\\\\{4b4bubF,ZwXa|bzuc0B/2/|b:kQoab;nOmxbGuKnb/ebabTpv,ebjbVrlrkylb?axxvb>bzb<a\\\\}b6z>uUa|3"));
$write("%s",("1bp5Q1aubp1bf1;nKx?aVbntq2bpm.Uakzu\\\\{Uahb.bdbwbcbb\\\\{1bZatxgrvb8.?l9*|vV*\\\\{b*sfb:d3b+/<afb4b<a?z2b\\\\{bIs+w0bCxF/7lD2Ra\\\\{,hbNa1bybtbQa+0,bZaJiXa7r+nfb@aybSz*elr7bvb9sfbaqjbwbmbvbFa2bVaQpEan3>a3l.2Z20btb=aibSrLs*b+/Ba.bPabbTzMyj\\\\}xf6+kbhbVaBqub7btq=a4bVr0+.+/+r\\\\{td\\\\}0zb>aOa2bu,lb/bayFaA,Oxr+>aar@a0bY*sn+bq0fljbMu\\\\}x<as.Tm3/6b3bBak-=aubXbu+Yr1bUadbrm;r;meuynE33b2yOlA,zbHl/k\\\\{bbbvbMwcbPaX\\\\}5brlOa--1b=aUqn,Iucb*wj|p|eb9*eb\\\\{bmbj|6mDaPaQa5blbFatb,,3b2z.b?q1b5bPaCa3b|*8rtbdw2q6,hr\\\\{bNalhhbFa>a4bIp.b;nNrYab\\\\{3bz+vq+exb0*W0ppNa5thb:kMrvlabWm>kabYa9y+xL*Wr|bQaj2J\\\\{E*\\\\}b@atb4|U|vbKx1bwbt1<xq2qyibnft1r1zb\\\\}bdwbwrpP,xfTqibbv8zSa6\\\\{,b*zxf0tQo*\\\\}0qxfXxOk/bV.5tNadb/b7bfbnrS|C|s.0b*b\\\\{b5bn1xbHsRpxf4saq|zdb\\\\{b2qS+j-WacbP-dx\\\\{b9bSaabkb7sbnFa2\\\\}tnjbz,MlO"));
$write("%s",("p;n6d6.Ta4b0b9*\\\\}cRpcb/bab9sNaSa5bfbu,s,myc/:0XaByQpdb.bOad.HrkyDl6b6bk,cwubbpYq4b=oix5bwbm,:mS\\\\{Caj.|b<xwbibLfGa.y\\\\{0Jd\\\\}mOa-bDoNa2xzbOa0b5\\\\{r|Na0k.b6bTa3b|0kbMnCp8ulbSz.b@aUaZ/vb-b>a+bTkChxvFa0bu-@yXe+b\\\\}b9kLpZasq\\\\}/vsnqFaXaBac++bVaPaT+0*6g>abwfnhbwq9rebCrxbdb6o0o2gp|Ta0bYaFacb.bTaXvCaTa\\\\}bBaumHzwb6wmblb0bXaEafb1b<wBaj.S+cbEs1qVa<vWaQaybp/nv;n|bcbpqyoSw<tkn=n9*|q5bDm\\\\}bJ\\\\{*\\\\}AmbbzbRa@w?o|bAovbkbtoSaRaFaAsyb3b8bEa3y|bWaubab|+Cae*Pa/bub2gtbabavlbSyWjCm@a,bhbgb2b>mubAa<hRqSkbb7babxfAwAayb6\\\\}DaXz,b>a/bzb+bXaRa*l|lu*5e=aCaGac|-bWaAalxAa.bYvVa\\\\{bZx?vCxMs*lB|Za4bX\\\\{8b/b\\\\{bEaCqybgbbbibwbYaUa|v1bD\\\\}xftbUakuSa?aXaxo8bB|k-=jVaeb9bZaCaAaJv3pkxgb>alhRal-9yirZaWpFaxb*bjbFaOk=wvxIxVw7,8bGz5bhbabgbodklubOadb2*vbBpjbJig\\\\{Sa0bFaQaMktb|b:s|+9*FaabyoabWvL|"));
$write("%s",("Ea5bZk,lDldbtbh+ibwqAafjCqRahbRaJi-m5b,bOxx|ab:zi,Tn4zBoq\\\\{cb5bZa6gBa=qzsdb\\\\}b5bdblbQa,q3p/b6bbbOaeb7z8ba|Y\\\\{Xahb=xabjbEmW*Da<kGnNacbbb\\\\}bXsPab\\\\{tbUyRatb:kTawblbbs=a*babVaXaDazb/b>a7r+knt\\\\{uxfQaKlFo-zzbrpol7b0bMv7bbzlbWpXaQaMdgbib6b0q>kjb=a|bib=\\\\}6\\\\{ir@sfv7bZajs<aubSa.qWa?aOa?o-bfb|bpyDa8bCe9b\\\\{b.byz|qHsavwbzb\\\\{dhb9kLrdx\\\\{f3bDsF\\\\{z\\\\}\\\\}s>nebNaCrMddb4a*|xfybFaRi5u7bPaWrYahfbbZt*zU\\\\}:wkbBxjb0kV\\\\}r*Q\\\\}|vSaTaEaS\\\\}=w9wa*VaY\\\\}hv8b9lSad*j|=aEa/bSaQaDeU\\\\}2bjbN\\\\}>rEaabWaTa@a3b:qAt@a<wOaRy>v=wPaWa@aSaEa=azbym/bTafb.kPailerdb6b9bEqCqbbybJ\\\\{6\\\\{XaP\\\\{<ecbUrAafzabP\\\\{vbOabqvtfq,tkzjb+bGaXp8b7s4|ct:wFa0o\\\\}b=a1q9v@angab|q/bAabqNax|Xam|1bYa6bbphbhbLuubbwcbUa>atbGaLlaowbkb6bBaebdqEaDa<ambxpYmzwl\\\\{mxib<a5bq\\\\{|\\\\{z\\\\{x\\\\{v\\\\{t\\\\{tiYyZatpxbNy\\\\{bwbn|1"));
$write("%s",("bmx5bNa0b;nxb-qzb5bubTaUakpolAzXaubAglb7s8bmb/bVa0rUg\\\\{nZaBaz\\\\{tbAg|zCavdsl/l3b8r:swbGamlEx4bHpCt3bJwabTa+bw\\\\{/bYq0q|vDawb2\\\\{Za*b>albmb:sDa8wcbup4x<aRaEa,bcbDambibfbZacbgbFp<a*w:p7!![2aba!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"g3b[2lpa\\\\})3(f\\\\{#(tnirP;)23&Z0bmbTaayQacbXn<acggbUa+b7bzb\\\\{babwb/bUaNaibafhbib+bzswbRaJpEawbBphbNtzbzbXatq?zjbQpNaCpPaPaebUa-btbup0bkuUaqdYajrdbup,b=a/bxhSaWpEaFacr6b*bfxHpWv0ytdstgbOo.bXaZaebxb4bmiVaEq/bftZaUeHj.wTaOkwd|bEnVaTaCaWalbRa>azoXa7blb>ais@ajb-bWmbbQl+b|kdb<adbcr5b2bFohb@a*bvtZavb4bRaoo/bFlYxsy|bSmoyjbWa5bkyhb6bYxvbYauslb2bFaibWaXxzbZakbDmWmfb/bBaMt8c-b=aybZa6w,bLq\\\\{b4beblbUaEaDeWaUa\\\\{b/bWambzbWaBa"));
$write("%s",("bbEa4b\\\\{shfCrAa>aUagb=aFaVa2p8rgbSa8qVa3bQovtRaDaubWa|g5bBa9v+b|vubbvEaGuOaupVakfcbwkAaebSumbxfibSaufvbEa6bebRq|bkbsoCaeb2bSa1bfb7b/bhtDa3b/b.tMufb\\\\{fxb\\\\{bngEaxfDaEaxbknAa@aWa=aSa.bRacbXrNaYaSk\\\\}uNo1s4aDjUt*bwb\\\\{b\\\\{b-o5bmbabGa=tDs;nOs?arvpqWa\\\\{uQaovSkBhGaMpQa0b?a:pibgbab\\\\{bkuXl8btbPazbDmfb6b2bmvng3bdb|beb=aWa\\\\}b*b>rbgyt3bhbcb>mdbBamb|bNa-bZsdb1bjq7bWk4bcl/obu1s*bjvYcdb6d<u+hYagbQa\\\\{bTaTaPaxb?acbElCa8u6b-bkb.bftWu9l1bQaFadotb/bEabbQaxpdb2b7b5n8bTa1bkbAm|k3bSa?s|bUaYaabmbbu2bul7kibtbGo\\\\{b*bXacb2bffQa8b1pqn>akb4f6bDa-bgbBn*b0bibdoQa3bDacb\\\\{bib1bar<aNarqCa+q2dabZaAa3bCauqwbUaisThFa,bib0bRaNayb*n4a4oyr2q0q.qqdPaNaBaxf6gJn|n?s-mzsZa/blbgbdombPaGqxfcb*b9bOnjb>a3q8bAa,bab*l9s9btbtb*kzb?a1bTkBa6b4bxf*b\\\\{s3b|sNaZaQaprHmXaXaOazb>s3b,bfb6q0bOp2b1bTaeb|bd"));
$write("%s",("r1bdbdoTaxbkb7mNp.bwb4bXakbPoWajbzbBa;n*b/b/s@azbubgb7bbpfb=ntbgb1sBaAajb0b4bym7bwbgb*bLqNa\\\\{blbvbXalbPa0bzbVa|b,bNavb<ajl8bhp0b|babBaFa*b3bnlFaYrwb*b+b,bOaAakbTaab0b,bXaEl<rGa\\\\}dtbBaUa@aYasm@a0kBbcbRpmb3bxbjnKoVa9pubxfBhXaTavbvbAa?b9bRa4nEaRa|bbb=aNaabPa8bvb=l2ogb4bdbiqvbDmyb*bmbtbdbkbOaJpYaRaAa*bmnWaabybQa6b>i/b+q\\\\}b;pabcbmmzbPaFa4b;n2bYafbMlEadb-buqabvbDaFazb3pCadb-lqdubUaub\\\\}b8b+bOaybkbWatbbbjb7bXajbgbPaXabb0bxbxbgbkbmbBacbab?aYavbNa/b=jzbeb1bcbjblhabibhbYabb\\\\{b+bxf8bZa0bkbSaOatbyb:p\\\\{bxfebvb2ncb\\\\}bOaBatb5kVakbgb,b\\\\{bgb\\\\{beb+bab\\\\}bSaSaHk/b2bPa|b6bkbFa?a/bgpOaTabbab>axfnmTk0b2dbpcb?a3bTaQlwbbbfbUaib,bPm.b-bRawb0bAo3b0bub>mNkfbwb7b8bTh\\\\}bTaZatb8b,bFawb.bCafoxokbvb6bjb0nubfbzb@aBaGaJmmoXaEe+bQaDatiriFj=lYaeb.bMfubrmWa6kOaiblbybDalbwbBh5k5b/bNm"));
$write("%s",("ynCaxffndnSaFk3b\"\"),\"& VbLf &\"(\"\"Wa7mdmxbabQaUa/bZa=ambmbXafbtb0b0bGaVkXaUaOa,bvbjbcbxlTaNa5b3bWkdnYa8b|nvl8babXaablbangb-f>aebtbTaub1bImYajb9b.b?aebzbNaCaBmRaXaxbQabb3bkb5bQa1bXamb\\\\{bSkcb8b2bfb-b+bfbQaAambbb8b9bzbjbRazb2blb1bebmb2bQa7b7ixf-b\\\\{b8b4b5bOaCa5b7bVaKlNa\\\\}bkbwm<aUa?aPaibTadbmb/m\\\\}bFahb,bdbRa\\\\}bxm>kdbQaub\\\\{bkbBa|bDaUaPa7bDa@aFa1bWa>aFa9bxb<aFa+bWa?kOaHf,kjbTa.bhb*bBaDafbJhcbmbhbvblbxfBa+bAklbYaZa-bib2bXaHk7bcbxb4a;lEjGj3b>ajbDaBaOaDakb=ajbubub*bAaFambEazbdbVbjbPa,bCezbmbSaXaFa6babzbxfmb,bCaFa-b7bTaQahb<aCa6bwb6bmbTkxf\\\\}b6b,bkbjbibvbVatb*b,bebBgvb@a\\\\{b-bhbaf.bjbhbjb|blbhb>axbzbEaubxb7bdbCaEaybLeQa4bSa>aDa*bibBadb9b*b-bEa7b6bAaEa:ifkzjckLjnjdjvihjYi8j;atjZi?aXitj\\\\{j8j-b:isjCa8jwb\\\\}c:i2j6iMjEa+i|jRi8jMi4asiCj9atiSfqi/b-b4b-a8guboftj+joj0j"));
$write("%s",("*i9aEaOatj-i+imjue:a-bhj=aAanjqj,inj4icj@a<aydTigjejhj>i-a<iWifj:aCa8aaj>aAa5i:iBc1iGiAaAe5iOijiwi@i8iBa*c;iCi*bLdqg,e5bxb|i9i7i5iwi3iOa|i/iBcAa*c\\\\{b\\\\}i0i.iFa@a-a*i|izi9awi\\\\{ixb8aCa@a*c*e8aviHa8arb8a8a2b4a4a3aRf4aNd3bWb6bfdzbxbubjcLfMfKf5a,d-a\\\\{d1bGb1bQgLheh?a=aRfJgjf4hhcXg=gVg>aBaKg|b|bvbag.b3bze?a3hfhMgBa?a3aHbXb8grbIgefbePgWdNgDaAeKg2b3bNf,gid:d-aue-b3aCe3aKa\\\\{b;aqdwbhfIa3b1b2g,b|b0atfWg;gCaKg.b,fefCdWfUfSf@aKgybIgtf<fXd<gBaRf5a3b9f1aCd1adcHcubwbxf,btfVfzfTf@a3a1bhfwb+b-aYbhd/b8bifXc;a:b6a5a-b;dZapghd5btgEf3bye7d5dNf-awb-f3b|d;a<b:b3b-a8b5d,bxb2b2btb;aefWd=fPa;f3a>a3alc-aLf/b3b4b.bHa8byb2bpdtbyexb5b+bAbefXdyf\\\\{fce9cteHa6f5eGawfxb-b6d4a-a.b\\\\{bndMaja-bPaBabesfGa+b,e?adfGa5a5a4d2bzb;azb-bWb3b2b5c?a?ace-aRaYaOaVafbVaibNa=ace?a;a>a-aVaNaUaievbpbEaed7"));
$write("%s",("bEaAaCa?a>anb,eubFbzbzeMa?dke<bFaFa9a>a:b;aocGd+b+btb\\\\{bvb3b:dJa2b-abdocZbXbVb;aie6azcdecejegeoc/abeRbZd6a/aXdbeXdIcUdRbWdCdBd9a2b5aMdKdIdGdxbvbtb+b/bxb1b5a1a/aCdhcockc/aFc:aIaXbtb,b:avb|b+bub4bcb-bqdodmdHaebdbJaGaxb,btb-b8a1bxbwbtbxbUa?b|b3bvbxbfbocnb5aXb.b+cXb-avb*c|c6awb-bxb6apbCc7bGa7bnbIcyc*b*bIcwc/adcgcRbccac>a8a?a2a6a\\\\}bKaKa6avb5aYbVa5aJa7bHa=aGa>a:aGaCaJa\\\\}b-a1b.bybjcoc|boc7aEaqboc2bsbsb/ahcbc5anbHa6aRbdcsb*bRbobQbNaHa3b-b|b1b/bJaNa/aob5a/a5a9a4a2b2a4a5azb.b+b;axb+b.b2b-b.bvb!![2aba!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"g3b[2lpa\\\\})3(f\\\\{#(tnirP;)23&*3~ia6(f\\\\{#,43.3\\\\}ea1150Y3\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'X4.ca06b4[b4[b4Soa678(f\\\\{#=s,y=z,p"));
$write("%s",("8Lfa59612j6[b4[b4[b4Nfa97571\\\\{=Pea5392Y3\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'d6[b4[b4[j8(&a3362(f\\\\{#=y,]99999[gnirtS wen=][c n3aea\\\\{)v]y3b&a(niam diov citats cilbup\\\\{RQ ssalcY8Mca75R6[b4[vBTpa(f\\\\{# cdln\\\\})0089#AUca17a4a/a;maertStnirP/oi/avajL tuo/metsyS/gnal/avaj[8bkategn\\\\})8027jCV\\\\}a655(f\\\\{#2 kcats timil.n\\\\})0294f6Vna587(f\\\\{#]; V);N;aM5ecaL[Z;aU;hpa dohtem.n\\\\})6332D4Uja53401(f\\\\{#K7noa repus.n\\\\})25992BUda9185CacaRQL5cgassalc.E>Lca76CE)C=/va251(f\\\\{#(=:s;0=:c=:i;)\\\\{8ajaerudecorp~5Lda970\\\\{4a~5Pda703\\\\}5apatnirp.biL.oken\\\\{$5bianoitcnufDC[$<dta918(f\\\\{#(rtStup=niamXONca04A5el:Mwa402(f\\\\{#(egnar=:n,i rof2@%n403a<0Z0Z/512152353/2/2166263=4/3141625>>914151:1/>5Ufat+)6,45Uea1312h5Xka(taepeR.S+n5Vfa41310n5Vda=:s7=c.acnuf;\\\\}r nruter;\\\\}\\\\})84-)n(tni,]1+2%%i:2%%i[74Lb"));
$write("%s",("a3\\\\}FUca7275acawW76VD8bja=+r\\\\{esle\\\\}o4TbavY3Toa=+r\\\\{84<n fi\\\\{s O?jz4Tx5Uka:r\\\\{gnirts)f3aea s(tm;a&=Ubaso4ad4TbaS|7Udatmf[3TjaF(tropmi;\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'Lafagakca7GMca32$Qa;Hax6Md4cba-Y3Tiatnirp te~9Mja115(f\\\\{#(nFKQca55qAa#a,s(llAetirW;)(resUtxeTtuptuO=:C;N&Ua*6ab4SdaS C[3M.3aca&(Y4Sba b6[b6TiaRQ margog5O.3ajaS D : ; Rm5Tba\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'X3Sqa. EPYT B C : ; Aj5Tka)*,*(ETIRWt5UhaA B : ;e4Sba [2cj5Vba:a4(+3[+3wda(nfOC&ba1lSa|aetirwf:oin\\\\})61(f\\\\{#>-)_(niamq3dvD~Q?afacnirpU@~na7(f\\\\{#(stup.OIhU,kWa|aM diov\\\\{noitacilppA:RQ ssalcWV~%JfR3diaohtem06x13kz6a.Xcpadiov;oidts.dts #Lay4\\\\{kaenil-etirwt6lva(,\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'s%\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'(gol.elosnoc;)\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'K3s[2cya\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\' nioj.)1+n(yarrA>-)n(=ff4kia!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\}54,1\\\\{.n3cja# qes-er(3Rdba&l5rba!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"URk$3lo3r33tla1% ecalper.S4l(3cU=gsarts(# pam(]YALPSIDq6cua!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\".NOISIVID ERUDECORPU3kma.RQ .DI-MARG~3oE3dnaNOITACIFITNED+:dsa[tac-yzal(s[qesod(n6apa!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\"\"\\\\\\\\\\\"\");\\\\}\\\\}!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\");\\\\}/****/e3a\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"),s[99999],*q=s;int main()\\\\{int n,m;for(;*p;)\\\\{n=(*p-5)%92+(p[1]-5)%92*87;p+=2;if(n>3999)for(m=(*p++-5)%92+6;m--;q++)*q=q[4000-n];else for(;n--;)*q++=*p++;\\\\}puts(s);return 0;\\\\}\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\");gsub(/!/,\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\",s);for(print\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"define void f(n)\\\\{\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"00g,\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";for(m=1;m<256;m*=2)\\\\{\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\"));
$write("%s",("\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"00g,4,:\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";if(n/m%2)\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"4+\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\",\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";\\\\};\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"4,:,\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\}\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"389**6+44*6+00p45*,\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";++j<=length(s);print\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"f(\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"n\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\");\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\")for(n=9;substr(s,j,1)!=sprintf(\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"%c\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\",++n););s=\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"4,:,\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";split(\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"145 160 17 17 17 23 252 141 0 46 125 231 229 231 250 151 243 243 243 231 231 207 159 63 4 231 249 255 191 225 17 127 206 103 51 57 152 37 255 57 204 230 103 48 79 159 159 151 252 231 51 51 57 193 47 249 204 230 102 115 4 251 190 249 243 207 57 206 115 158 9 231 57 156 206 102 9 193 48 96 22 236\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\",a);for(i in a)\\\\{s=s 0;for(c=a"));
$write("%s",("[i]+0;c;c--)s=s\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"1+\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";s=s\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\",\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";\\\\}print s\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"@\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\nquit\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\}\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\")');\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";FORiTO UPBtDO INTn:=ABSt[i];print(REPR(50+n%64)+c+REPR(50+n%8MOD8)+c+REPR(50+nMOD8)+b+\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"J\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"+a)OD\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\"\");end;\\\"\")\\nsys.exit 0}\"\")]]></xsl:template></xsl:stylesheet>\":s=\"   \":For i=0To 7:s &=Chr(32-(Asc(c)>>7-i And 1)*23):Next:System.Console.Write(s &n &Chr(9)&n &\"  \"):Next:System.Console.Write(n &n &n):End Sub:End Module"));
end endmodule