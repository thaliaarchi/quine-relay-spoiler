module QR;initial begin $write("%s",("let s=(\"Module QR:Sub Main():Dim s,n,i,c As Object:n=Chr(10):For Each c in\\\"<?xml version='1.0'?><?xml-stylesheet type='text/xsl'href='QR.xslt'?><xsl:stylesheet version='1.0' xmlns:xsl='http://www.w3.org/1999/XSL/Transform'><xsl:output method='text'/><xsl:template match='/'><![CDATA[sub f(s$,n)print(s$);:for i=1to n print(\\\"\\\"\\\\\\\\\\\"\\\");:next:end sub:f(\\\"\\\"write,format=\\\\\\\"\\\"%s%s%s%s%s\\\\\\\"\\\",\\\\n(\\\\\\\"\\\"\\\"\\\",2):f(\\\"\\\"write{-}{txt}{echo -E $'(\\\"\\\",1):f(\\\"\\\"\\\\\\\"\\\"with Ada.Text_Io;procedure qr is begin Ada.Text_Io.Put(\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"interp:library\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"afnix-sio\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans O(n)\\\"\\\",2):f(\\\"\\\"{trans o(afnix:sio:OutputTe"));
$write("%s",("rm)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"o:write(Byte(+ 128 n))\\\"\\\",2):f(\\\"\\\"}\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans f(v n)\\\"\\\",2):f(\\\"\\\"{\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"O(+(/ n 64)107)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"O(n:mod 64)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"O v\\\"\\\",2):f(\\\"\\\"}\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans D(n)\\\"\\\",2):f(\\\"\\\"{if(< n 4)\\\"\\\",2):f(\\\"\\\"{f(+(* 6 n)9)48\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{if(n:odd-p)\\\"\\\",2):f(\\\"\\\"{D(- n 3)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 27 48\\\"\\\",9):f"));
$write("%s",("(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 36 11\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{D(/ n 2)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 21 48\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 48 20\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans S\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"STRINGz:=REPR226+REPR153,a:=z+REPR166,b:=a+\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"2\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"+z+REPR160,c:=b+\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"8\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"+z+REPR165,t:=\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"#include<iostream>\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\""));
$write("%s",("\\\"\\\\\\\"\\\"+REPR(10)+\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"int\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"+REPR(32)+\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"main()\\\"\\\",2):f(\\\"\\\"{puts(\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"class QR\\\"\\\",2):f(\\\"\\\"{public static void main(String[]v)\\\"\\\",2):f(\\\"\\\"{System.out.print((\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"write(\\\"\\\",4):f(\\\"\\\"'implement main0()=print(^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"BEGIN\\\"\\\",2):f(\\\"\\\"{print(^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"echo ^\\\"\\\",4):f(\\\"\\\"'f(s)\\\"\\\",2):f(\\\"\\\"{System.out.print(s);\\\"\\\",2):f(\\\"\\\"}s=^^^^^^^\\\"\\\",1"));
$write("%s",("21):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"389**6+44*6+00p45*,^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";for(c:(^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"#include<stdio.h>^^^^^^^^nchar*p=(^^^^^^^^^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"Ra#include<iostream>^^^^^^^^^^^^^^^^nint main()\\\"\\\",2):f(\\\"\\\"{std::cout<<(^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"class Program\\\"\\\",2):f(\\\"\\\"{public static void M83abbSystem.Console.Write(^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\""));
$write("%s",("\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"Quine Relay Coffee.^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^n^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^nIngredients.^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^n^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");for(int i=9;i++<126;)[3pva$^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",2):f(\\\"\\\"{i\\\"\\\",2):f(\\\"\\\"} g caffeine \\\"\\\",2):f(\\\"\\\"{i\\\"\\\",2):f(\\\"\\\"}I3b54rja^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^nMethodv4f#ae"));
$write("%s",("ach(char c in(^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")))^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^[2al3dp3c[2cs3c,3l[2k@3kqa^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")s rts(ec"));
$write("%s",("alper.h3eja^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"     53c4a SUTATS(egassem^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"rts(nltnirp(])]^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\".NUR POTSu4cba.C3dh3dX3bba[65bX4df5lp3lna\\\"\\\",2):f(\\\"\\\"})1(f\\\"\\\",2):f(\\\"\\\"{#\\\"\\\",2):"));
$write("%s",("f(\\\"\\\"};)06xt3dba;+3noa3(f\\\"\\\",2):f(\\\"\\\"{#qp]\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"};)0,#3rv3rR3sv3mba723284-fa(f;)1q5.ba.>4[ga#(f;)3P6[=43ba7=4.<4[<4[<4[v3gJ=d=4[73++>u?4[73xda,43?4[?43ma^\\\"\\\",4):f(\\\"\\\"'^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^\\\"\\\",4):f(\\\"\\\"'^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^\\\"\\\",4):f(\\\"\\\"' D ; EYB RCo8[.6[?4;ba5qB/daDNE&6[&6[&6[8Emca AL9[)6[)6[v3oeaPOTS^\\\"\\\",4):f(\\\"\\\"'^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^\\\"\\\",4):f(\\\"\\\"'^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^\\\"\\\",4):f(\\\"\\\"'6[^\\\"\\\",4):f(\\\"\\\"'^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\""));
$write("%s",("\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^\\\"\\\",4):f(\\\"\\\"'^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^\\\"\\\",4):f(\\\"\\\"'6[^\\\"\\\",4):f(\\\"\\\"'^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^\\\"\\\",4):f(\\\"\\\"'^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^\\\"\\\",4):f(\\\"\\\"'6[M9pL9[(6[(6[v3moaRQ margorp dne16[16[16[v3lbaST9[&6[&6[JQ[~6[?4Nba4~6[~6[~6[~6>ba&g=[$6[$6[.@neaPOOL|N[,6[4@[>Xp>4[#6[#6[#6[#6[?4Kba4yGXk4dba0j4[fa#(f;)980da&,)&?[=8[b<[\\\"\\\",2):f(\\\"\\\"{Wnga. TNUOOB[,6[,6[83nearahcGI[)6[)6[R9ogaB OD 0~W[-6[-6[;Po33)$6[$6[;PBca)Av=[&6[&6[cToYS[^\\\"\\\",4):f(\\\"\\\"'^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9)"));
$write("%s",(":f(\\\"\\\"\\\\\\\"\\\"^\\\"\\\",4):f(\\\"\\\"'^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^\\\"\\\",4):f(\\\"\\\"'6[p=[v3nqaEUNITNOC      0136[36[36[sDnV9[&6[&6[lDoG@[^\\\"\\\",4):f(\\\"\\\"'^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^\\\"\\\",4):f(\\\"\\\"'^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^\\\"\\\",4):f(\\\"\\\"'6[^\\\"\\\",4):f(\\\"\\\"'^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^\\\"\\\",4):f(\\\"\\\"'^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^\\\"\\\",4):f(\\\"\\\"'6[G@sba.)6[)6[)6[@4mja1=I 01 OD-6[-6[-6[C@neaA PU*6[*6[*6[v3mxa;TIUQ;)s(maertSesolC;))T4[96[FN[v3kfatiuqnp41ca46p4.N5[3"));
$write("%s",("7[?4:ca11o;/072ca82m4/g<[27[?4;da932A4.maetalpmetdne.>72ca65y4/>7[>7[%D<ba9G@/ca\\\"\\\",2):f(\\\"\\\"};&6[&6[f;<ba1JG0ba^\\\"\\\",4):f(\\\"\\\"'^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^\\\"\\\",4):f(\\\"\\\"'^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^\\\"\\\",4):f(\\\"\\\"'@4[%6[oK[#6[#6[#6[#6\\\"\\\",2):f(\\\"\\\"}damifo=[(6[?4<ca37WC/l41ba0j4[)Oada923g<[=8[=8[+?[#6[#6[#6Qbat?4[$6[rV;ba6ZL/^\\\"\\\",4):f(\\\"\\\"'^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^\\\"\\\",4):f(\\\"\\\"'^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^\\\"\\\",4):f(\\\"\\\"'?[j47da601^\\\"\\\",4):f(\\\"\\\"'^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):"));
$write("%s",("f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^\\\"\\\",4):f(\\\"\\\"'^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^\\\"\\\",4):f(\\\"\\\"'?/%a315133A71/129@31916G21661421553/|7[a9[&<;ca76Q7[a9[j4fda298BG/ra%%%%\\\"\\\",2):f(\\\"\\\"}*+1%%%%811 -$:2ca19/5[:6[j4gba8<<0haj:+1 j@>:[#<[?4:ca62#<[C8[=Dhca49#</bawX6[=8[dH;ca7827[=8[U:gca96EVX<8[<8[?4nca11iQ/=8[j48ca54=8/baWY6[>8[?4:da263>8[>8[<Ohca02>8/ba\\\"\\\",2):f(\\\"\\\"{Y6[>8[?4;ca06>8[>8[j4hca69x5/bann41da468+6[+6[(>hba3k<0):[j<[kM;ca85=8[=8[IAhca283X/x5[j47ca75V:0wa)(esolc.z;)][etyb sa)^\\\"\\\",4):f(\\\"\\\"'^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^\\\"\\\",4):f(\\\"\\\"'^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^\\\"\\\",4):"));
$write("%s",("f(\\\"\\\"'09[q;[?4:o;0#6[#6[#6[#6mfa2200uq42ca84G?[.=[G?[x5[x5[x5[x5[x5[x5[x5[x5[x5[x5[m4[x5[x5[x5[x5[x5[x5[x5[x5[x5[x5Gba2EP[EP[EP[jT[#6[#6[#6Rba,%6[%6[%6[E9[#6[#6[#6~ba!m41ba6m4/ca~~37[37[37[S:[#6[#6[#6~ea(rt.(6[(6[(6[H9[#6[#6[#6~ba)BA[v3cda\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"};p4[SBfdadnes4[s4gra~~~~PUEVIGESAELPnr3ala~~1,TUODAERw3a:4[:4i$a(etirw;\\\"\\\",2):f(\\\"\\\"};u=:c;))652%%%%)u-c((||54[54ida#-<u4[u4ida||i15[15lhaBUS1,ODz4[^\\\"\\\",4):f(\\\"\\\"'^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^\\\"\\\",4):f(\\\"\\\"'^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^\\\"\\\",4):f(\\\"\\\"'8pka)3/4%%%%i(g:c4;[04jr;[r;wPa2=:/t;2%%%%t+2*u=:u\\\"\\\",2):f(\\\"\\\"{od7 ot0 yreve;i-=:u;1=:+i\\\"\\\",2):f(\\\"\\\"{od))1(evom(dr"));
$write("%s",("o=:t elihw?s;)s*z9[L;ny9[y9uz4[z4i0Adladohtem dne.s3dganrutern3dCaV);gnirtS/gnal/avajL(nltnirp/maertStnirP/oi/avaj lautrivekovniJ3d25[25i[2cib\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"};0=q;)]q[c=z(tnirp.tuo.metsyS;)0(tArahc.y+z=]++n[c;y:]q[c?n<q=y\\\"\\\",2):f(\\\"\\\"{)0>2%%%%++i(fi;48%%%%)31-)i>3c&as(+87*q=q\\\"\\\",2):f(\\\"\\\"{);01902<i;(rof;n)rahc(+O5[O5q[2k.4[.4%oa=]n[c);621<n++z6aqa0=q,0=n,0=i tni;R4[R4%mc6aVh4asdRbQeKkxfvfDk8f<bedRbkkP=;agb-a|dzdxd8fGb8aqeRdYd5amF\\\"\\\",2):f(\\\"\\\"}i;agb-epb>aqeRdHa>aJaRaAdteFbae:b6aOa5aachgXzN\\\"\\\",2):f(\\\"\\\"{9aV\\\"\\\",2):f(\\\"\\\"}4aLa7a;a4a<a2hGlkdxd;aNa?c6a|eebHaFaIaebzeJaeb9a\\\\\\\"\\\"),\\\\n(\\\\\\\"\\\"/a6a2dQbUe-f2a-f9aV\\\"\\\",2):f(\\\"\\\"}5d6cRbC3g3c-f/aof0f8fHg5a+h5e,V2e6aRa;d0rMfi*\\\"\\\",2):f(\\\"\\\"}h;aTapc4aLcEeVhof6amcylsbRg*\\\"\\\""));
$write("%s",(",2):f(\\\"\\\"{=fybxcxc@:UeAa2a6aZf7a6a@a1a:a?aMbKaKa6a?e:as,2a?a@fMbAfGa>a:bXfEl;f\\\"\\\",2):f(\\\"\\\"{bHa4atc\\\"\\\",2):f(\\\"\\\"{iNauEZsX\\\"\\\",2):f(\\\"\\\"{Zs\\\"\\\",2):f(\\\"\\\"}bJaMa\\\"\\\",2):f(\\\"\\\"}bJaHz/9JaJav;JaMdJa8b;w;a51TaKa51Ta8bm?kCPalPN69EKa8bN6?aTa51\\\"\\\",2):f(\\\"\\\"}3aqalC=sJaLaJa8b2-Naf4cya8blC4blC:bZsuEZsuEkCJaHay3aca=sk3a)aFd7=;a8b|t:aUa:a;wRh9f7f-l4a?6sbsb2be3^\\\"\\\",4):f(\\\"\\\"'^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^\\\"\\\",4):f(\\\"\\\"'^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^\\\"\\\",4):f(\\\"\\\"'maRhDa-a|bY\\\"\\\",2):f(\\\"\\\"}-a46asaa*Ue>ajj1aKaKa?a@ft6cga2jobdgx6csasbRg*b-a/bxcHa|fQ-e3c,c\\\"\\\",2):f(\\\"\\\"}b1aMg1aTfXf\\\"\\\",2):f(\\\"\\\"{bHaQ-8f-e:a:a\\\"\\\",2):f(\\\"\\\"}bHaYfJa\\\"\\\",2):f(\\\"\\\"}b5aAd"));
$write("%s",("te@aXfeiQ-xcpb7anb2b:b1a2fuj@d<f6aAjxcHa>aIfGfHj-a;fei-fHamcdg9f|fQ-ze6g-fHa<k;a/aah<bbhlh<apb/aahlhnb<a<a7b:b1a/aah/adgbgFaai|b1aGa3b:b1aphHaQ-HaUebiCe|bxc3b0a:b1aIa|bzeJa|c5b#aQb-f<b=a-atm*c3bxdUe=a-a?a,H9ai3edbAg7apbEQMgKgIgGg9apbNgLgJgHgKcdc/bPcgfvf1h,h7aEQokmkMatm*cEc,dJa>a2a:b6aUijkMa?a,Hri+c>h6a13idbxdtbfCng/aah=aLhRalbOaCdlbOaf@k+NaLh:k9h7b5a<k8fwbXiUe2b5aog:i4b-bhcEm1i1iAo0c/bxd;azbgiJiq?aea6a2b:>g5a\\\"\\\",2):f(\\\"\\\"{S6aan2a5aBm.;6aFjfvji9h7hAmHa1dmd.hHaZfmiAkHapbi3a2bkl<b3bxd6a+h\\\"\\\",2):f(\\\"\\\"{k2hfljbGhGhvftf\\\"\\\",2):f(\\\"\\\"{z;a,b1hq8fbpbubld1bZb5Q+iZpNiEc,dFj8kij<b<b<b\\\"\\\",2):f(\\\"\\\"{j:bqj<b<b,c,j\\\"\\\",2):f(\\\"\\\"}j7b-b,jEapn3bDdfk/i9a7blg-a5b@Y,c,j=a9a7bFtq3e13ecaxj13ceaEzikA3c/3ggaJb7bCf#3bxD1ba0wD.$ak9jAa>a6z9a9\\\"\\\",2):f(\\\"\\\"}xb-a5bh7UjKizk,c,ji3a)aD"));
$write("%s",("lNvCg,c,jsb8fFj8k8jyjCa.i6a3iljDjiji3aia@kdk<bze0DegaFj8krk-3crb,k*k3a6a<bGh>i-;2b2a2az9AjxkeiwbXi8f*3nc:e-bJaJaubph5a=f=anbAjybYj5a,bJa6a7b5a8gwbXiHa:e-b9a9b9aIgAjWf>am3awa@a@aAjWf*3:a|b9a0b9a*3-CaAa>e|b3g9bJa0bAjWf-b9aIg9aCaAaJa9bAjnbJa6a|b5a,b8f:e-b5a<mtb-aR<a&aVh,OwSRhz9Wf8bAd\\\"\\\",2):f(\\\"\\\"}h-az9*bV--az9Wf7s3h13a5aXb;d/g/bxd6a-b9a8b9a7bJcJaybim>aGh>aJa*c@dxc?brso3a1a-bxlteUe*3:.KdP6vb:atcJaub5aEcxb-4,b4b-b9g8f77aia6k3amd.ho3a#a@kd*.ipb;awbXiVkAm\\\"\\\",2):f(\\\"\\\"{S4G,O|Q/I.;F4aphFcClXk/mOmsl4lencnvmyn.mTlpl,OTZ,lA\\\"\\\",2):f(\\\"\\\"{Tr;xexVGJuQwGhn/,nzojb,nzo-bUj+ysLP1Za<qm-k9vb=/W;.vZa@niulbAqZalb|*\\\"\\\",2):f(\\\"\\\"}65QtIEwxo,nex@\\\"\\\",2):f(\\\"\\\"}gb<a>aZahb=atcuppqgJP?ub,YYa*UD5tFNoToFE<apqjbC=n.zzuvhGGv1r>av9Wak:FqjblEjvEC=atblbTa|bT0C?1,hb3bVYmb6Hy8tDtBopgbOar@v"));
$write("%s",("bZ|bbiu;p5bmbInVa*F@G\\\"\\\",2):f(\\\"\\\"}vTpYMX*ptJ9LBS,V5ybPtA>fo2skb6b.>89Eg/bkyou+|l?cUI-CCmb6b|b:u\\\"\\\",2):f(\\\"\\\"{dt29bxx*bybVh,OTZa18LUa+qDyC1R,/JZvFG+*dI,d\\\"\\\",2):f(\\\"\\\"}0tiYajYzpAa.h9/iKvbc4Ut6oq*<acbSxubdbU1\\\"\\\",2):f(\\\"\\\"{b6+KovoVaCazPA.*hYt;\\\"\\\",2):f(\\\"\\\"{QaDyjb6N;p+bn*Za\\\"\\\",2):f(\\\"\\\"{bSa/5U\\\"\\\",2):f(\\\"\\\"}.>|brs\\\"\\\",2):f(\\\"\\\"{PAwldU+O7wp:7TaP8U;\\\"\\\",2):f(\\\"\\\"}U:ncEnAp6*d9AEslCQ/01<am8>\\\"\\\",2):f(\\\"\\\"}3b@y9b7b=yEaPfI5>/qkb\\\"\\\",2):f(\\\"\\\"{8b7bMt?*n-s;h96Oi\\\"\\\",2):f(\\\"\\\"{Hp=rUHN1+bAqe1\\\"\\\",2):f(\\\"\\\"{7FaZ.NaLU3Oc\\\"\\\",2):f(\\\"\\\"}vyyr>wZIO*y:o9PMoPPix/TaAa/burU+DazLTaoAG>+3:9Mr:n|6a\\\"\\\",2):f(\\\"\\\"}d0RPf\\\"\\\",2):f(\\\"\\\"}v3+Rw,b,SWLGo6bh:OKAaYa\\\"\\\",2):f(\\\"\\\"}b4?Oax,AaYa<HIzir:9dbwb9P,Q9sQu\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"{l,f1*b>ahS|0f1=:CgNRCgNoh.@NZIp?bbrSJJ6bZH.P3+O"));
$write("%s",("y7J,oU06ylbDa|z3+fq+qePcPaPjp<DAa@akqEajb?aVulNMO-7=PS3J14SjbuBwPA.DalBmR=aC\\\"\\\",2):f(\\\"\\\"{jbDar\\\"\\\",2):f(\\\"\\\"{DamblbDavb97,bCze\\\"\\\",2):f(\\\"\\\"}<5|boNlbz6rwkQlb-oDaU=,p4bupF?=a*4U=,pzie=mbNa3+wr:nPimbNambUgsv,nXa535wdO\\\"\\\",2):f(\\\"\\\"{|.b,&6bpdeGR\\\"\\\",2):f(\\\"\\\"}uoz6GhuN3+4b|0||\\\"\\\",2):f(\\\"\\\"{rZalb=:q|K524,QqPk<=N,QQakbSaIn+|:nQP3+SiTaX1LZeG,QavOa3+iU:nvb7+AQ7z*nrN@noNlb7\\\"\\\",2):f(\\\"\\\"{f0jNhJgN|qsyML0R,byb;+CaF?=aev;+,p7b/CnBNoDaoDBanBNo;qtFNa;+ub;q5PgbCaI\\\"\\\",2):f(\\\"\\\"}Q/gJx+l7rp+hGU\\\"\\\",2):f(\\\"\\\"{p7b:pwukuYwV6UtAx*D=aro6p0M0b;\\\"\\\",2):f(\\\"\\\"{X|sr-MJJ.bHT:Gnrm+T;0BG>l?D*-bbp0<AaYaVI30Pn6Ln2pM-HHT1Qt6aqaTaTL?ajb2bB:ep?Yo3aza,bJJ5pdPEasr+b<a>nn2swno4%3dMcg1UH4p7bqkCw/b4poPHTZ.<aDa+b<a>aiM4pmb@GfbewTaPa*g:swwubtblL:sWYipeb2<jblB\\\"\\\",2):f(\\\"\\\"}bcb@atb4bcLtbaL9znw"));
$write("%s",("WK?5TKRKe+ToL?T0ZavW,yNEFKDKwbvWk\\\"\\\",2):f(\\\"\\\"}DaEaoDA=oDDDablUX;fbtbBabb<a=ajb0Q.-RCB.ExKPvb7bM.DyU5k.i\\\"\\\",2):f(\\\"\\\"{-bXu?8==*brka8HU*bDaHT,zr|r46nub|\\\"\\\",2):f(\\\"\\\"{3b;xM4bpAQ<aTa=yI4NJ/g/bVh.Dg\\\"\\\",2):f(\\\"\\\"{de5/bhbabTaesAqesebot\\\"\\\",2):f(\\\"\\\"{bkoeo1bH|-dZuv-AyXOVOTO|4domr5y5beoio?S5bhoeb<2xb:sO01:ghb4z6tbB,ZaSrCwmo\\\"\\\",2):f(\\\"\\\"{,G;TI\\\"\\\",2):f(\\\"\\\"}b>IRakb5soPgBLpA>ao=ar7@X\\\"\\\",2):f(\\\"\\\"{,G;p.Ca?S9U8qVantmr>Idp5sA<;Ylthb3b7TO?TamKc=cbe,Ml2wab|bqtJ3+Q\\\"\\\",2):f(\\\"\\\"{LcbQHL2V>m.b3U0f*lb7Vhb*F3b/bd58bbr1,Yuy+AaA<Vy8E9vOacb.bxbRazFoRPolR.TTwt63bUpHodbZK-NQa3,W\\\"\\\",2):f(\\\"\\\"}WAd,6jqd.=a5X9s\\\"\\\",2):f(\\\"\\\"}LBjbf*3Rb\\\"\\\",2):f(\\\"\\\"{Tan@=Gvb+bAU+LDzUq>@PK|bTaMO0bOaZ\\\"\\\",2):f(\\\"\\\"}zb@118quTaa0tvMReq?al?Ta1\\\"\\\",2):f(\\\"\\\"}dp-b:B@OtPzbF+bx|5uIFaI+-y+Q|uss.b@B6bJzBs"));
$write("%s",("mzRZ2U5FPaQMi|rui|ur>*IU@a?:C-\\\"\\\",2):f(\\\"\\\"{G;?Sr\\\"\\\",2):f(\\\"\\\"{Rgb.bw1f*+r|7zrWaK@RZCa5bjbtFS|cbP|XO>t/b2r1+5Qg|6;\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"{bEPB./ElrldAU1|JHq=+w51n5GaeOCQE/y4Zacb6r4b|-24L1Ual2M.OZ,bMZKZIZe\\\"\\\",2):f(\\\"\\\"{GbrdYaXa.Xsq/L7,G;5Ah3J7H7h?|z9S5>ivirn-*\\\"\\\",2):f(\\\"\\\"{aN\\\"\\\",2):f(\\\"\\\"{bdwKKGups5b*y4qQZZTzo/CZ\\\"\\\",2):f(\\\"\\\"}Aq6|3XwbqItb7b2JNazjTa1\\\"\\\",2):f(\\\"\\\"}R\\\"\\\",2):f(\\\"\\\"}G\\\"\\\",2):f(\\\"\\\"}ubtbH<jy\\\"\\\",2):f(\\\"\\\"}:-bf*=vP1Gvebyb<aUa7-2ry1l,7-+rVXpo9sy@5FQ1\\\"\\\",2):f(\\\"\\\"}b\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"{=97oU1+rR3\\\"\\\",2):f(\\\"\\\"{r9RvDzoU=UDrv;wX32x8|rqgb\\\"\\\",2):f(\\\"\\\"{rU1VaO\\\"\\\",2):f(\\\"\\\"}B\\\"\\\",2):f(\\\"\\\"{uLW\\\"\\\",2):f(\\\"\\\"}e8Z\\\"\\\",2):f(\\\"\\\"}|*?A-yh\\\"\\\",2):f(\\\"\\\"}+Je\\\"\\\",2):f(\\\"\\\"}<5tb5?RoM.|b<a4bLIZ\\\"\\\",2):f(\\\"\\\"}ZaWahbm?m+yUB+Cav"));
$write("%s",("b0bS1w2jOYa3\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{<Va<vg?Avwrv6a@bzPn\\\"\\\",2):f(\\\"\\\"}t*uyYx01<RTw6syuYaPV8uaqnB9J-tA<<aOy/E+,-oL-Wa0x-b-zWy9NZkzv\\\"\\\",2):f(\\\"\\\"{|+sdb:\\\"\\\",2):f(\\\"\\\"{d5-b.v+qj0-/*b5Me1;*0<sR.pH?0<XaxX-oh<HihGK57@yb?ab.lbSD5bFttbHiEaV0qAe+c+m3a8bW;utJoaGuBz2wW+yT0z<6swb@a20C2lbOZSjTOZqk\\\"\\\",2):f(\\\"\\\"}borK@a.><2Bvd+b+uv5/dbUa<aVa=aA=VacuxX3y4bxba-Pah?Ca1btb2b=aZIM+HP3ylb7qR*Va1bibesaLmb\\\"\\\",2):f(\\\"\\\"{,0by,e,9+&6a&d.b\\\"\\\",2):f(\\\"\\\"{;K:>a9+C?>VbMkS?aVs,w01?a*pQqdqJqQaQM-bYx01NaKr9M=h6bDUaPXaPfi*Cavb\\\"\\\",2):f(\\\"\\\"}bC?Ju3b/bhv*phJB./EzoL\\\"\\\",2):f(\\\"\\\"}o2@tbw,b*UMkDH?YBaEzqQ7bgU1btb62vbGpWanyTa|J;sJzvBs?zz,4/J,nc,aCSa|zU\\\"\\\",2):f(\\\"\\\"{OaVLuM-HnLvbj8abAuIzX2gBybevnvqA0:Pf?.PfkwVvU<cb>q=hVavv4bM+GtoBibJt5b7bM.o\\\"\\\",2):f(\\\"\\\"{kbQ*wbB0|-Dq>a7Vs646Ta7bUWbr.bB*@"));
$write("%s",("a4p*6G2\\\"\\\",2):f(\\\"\\\"}:cOjb\\\"\\\",2):f(\\\"\\\"{b:ss;Aq*6azdJ\\\"\\\",2):f(\\\"\\\"}0bq|c4@GeKZa*,lNWEsL2b:v|G<a<v+d1bk\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{b:s40EAorLrhbR9vbo3j-Gsi\\\"\\\",2):f(\\\"\\\"{<?imLxYoX@EakyZaZrOG>a=ar-c:U*Val|EDabXn7bib4+Xix-*vXzZ6BqmbY6vwZtub3,5zR/Q=w+,o;qGl,Qbb|J@KCa7b=aqiO=5Mkd6bM-+|J3=VFa|rTwSaotGh8:@XQQYahv\\\"\\\",2):f(\\\"\\\"{7zo-bSybxGyzoaU:uZ.hvPP-bSyc\\\"\\\",2):f(\\\"\\\"}pMs7uDe1bM+q:nGj.X;PQagtO*/\\\"\\\",2):f(\\\"\\\"{-brs5|lNt2lNQa*ztbs;ZNJz>a~6aqak5\\\"\\\",2):f(\\\"\\\"{rZa5bNa3n5>tb4BahaA5^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^[2fha\\\"\\\",2):f(\\\"\\\"})3(f\\\"\\\",2):f(\\\"\\\"{#v3r"));
$write("%s",("ga(f;)0,73-|bzv\\\"\\\",2):f(\\\"\\\"{bjbGQl2Y\\\"\\\",2):f(\\\"\\\"}evMr>sP-NSH\\\"\\\",2):f(\\\"\\\"{rp=aeb-b+JebsL\\\"\\\",2):f(\\\"\\\"}3a3|57bWNQo<2ti|RtiHMC=DMUDgqYaYn>awb,xb,F*J\\\"\\\",2):f(\\\"\\\"}PwsGlbHVKrfb-7U5dY3bVR=nqsF-Va-3cqabPkboDVRNaWqctUad4a(be,jxcsbb<H-bGhx2Q-Ts33VR2r\\\"\\\",2):f(\\\"\\\"}rjvpq;nGp*bUOC7F*DQh9NaAa@aNa*nlN>t\\\"\\\",2):f(\\\"\\\"},\\\"\\\",2):f(\\\"\\\"{n:->AtbWy6b0bOo2bCAr;gBWo:uWV@ae-T4\\\"\\\",2):f(\\\"\\\"{0Vawp6Olbzveb0girTwmzZDc5ablvbO\\\"\\\",2):f(\\\"\\\"}B\\\"\\\",2):f(\\\"\\\"{+*T|A36oZ@RaJ:PBwtPa?B.w;Zv,,bKAdP7zc0yb#Ca^\\\"\\\",4):f(\\\"\\\"'^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^\\\"\\\",4):f(\\\"\\\"'^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^\\\"\\\",4):f(\\\"\\\"'a@-<a>Pyb-xBvOp.>VpGQ3n.t0bnK5qusNS%3cDbNa9rDP7b;sWa"));
$write("%s",("?XQadq?<n5\\\"\\\",2):f(\\\"\\\"{4roQaQ>2sIHFas5YqmF\\\"\\\",2):f(\\\"\\\"{v3v;pkA=rEzmbR,<aQ7*bRa\\\"\\\",2):f(\\\"\\\"{|kdvAnw+Q+bXrAQ5qf0zbQp<aQE+Z*FhShbPa:\\\"\\\",2):f(\\\"\\\"{=:CqibPWSswb<rF,-wWOUOef61F-8\\\"\\\",2):f(\\\"\\\"}Vp=nNASwFAgpn*;3akaC?NacbpJquq3cmapoFt=:wq?S*/|6a^\\\"\\\",4):f(\\\"\\\"'^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^\\\"\\\",4):f(\\\"\\\"'^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^\\\"\\\",4):f(\\\"\\\"'cwbL3E\\\"\\\",2):f(\\\"\\\"{<uzbppb@o:5bNa8uuE,b4b=,=,mT9bAwPajyp?>pTAubVK.:8bhbh34wLu+4qk+2mRM3L6Qaf8V7O*CwS3lOivEfevs:Za4blbU+/b.b<qCwbQ2b6bfUCwAalbF|jO2blDov0D8r;w*b<ab47b|W,-|WktubBafwmb/yoDfUru<pNtCaZ\\\"\\\",2):f(\\\"\\\"}8TZa5bC?ebV\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{|b23n-|>tF|f:aVa\\\"\\\",2):f(\\\"\\\"{bXu1bgJ48"));
$write("%s",("lDQZTa+AC?j-QaO\\\"\\\",2):f(\\\"\\\"}<G6b-ydM/n/bibL3yuYaF/DaXaoVe?iAE-.0eGIJmdqWoV6AbbRaNSbIKb~byD?aoVabtv<gxTQZRnvDCavbRLjbGuRuoDV>yb3R8rOqq85t:Szjl7<WUH+v|blbrqccjbZ\\\"\\\",2):f(\\\"\\\"}=:/E+bLC:S;\\\"\\\",2):f(\\\"\\\"{GqTaGZy4ouVBoVZ6Na6I<vacO*+|KuvfH>(ba7d?vS?vba7S?.da,43?4[ha(f;)932A4.ia(ntnirpnt41da821t4.ba)T5[97[97[v3l2b<WY*W*V6LU+xgbZuw2wrvooDw2cb|-X14z7A1bjb;qp+wq\\\"\\\",2):f(\\\"\\\"{N:Sog.bmbubI>9wzo,4X:Xr\\\"\\\",2):f(\\\"\\\"{<<7CsKABvm22RQaFGF+hgYqWqlbBs2UsNz|NSXnrsUqZ0cr,-jbcRGvFa\\\"\\\",2):f(\\\"\\\"}b6wi3csaJ<8ySz8b;H6OecR:Is#Zisd|C\\\"\\\",2):f(\\\"\\\"{<hXyrM.OtMtybEsPtbtbbRodw>a;1s+9pCxF5Vadb\\\"\\\",2):f(\\\"\\\"}p|iG</bAaYaTz*n7@yba5BaK2cbdZ<alb+-cuEKQH3b-5+5\\\"\\\",2):f(\\\"\\\"}5\\\"\\\",2):f(\\\"\\\"}@.8,2v5b;P-bbtHQFgyubFXqtxbQaZRYa4+,|*v-6ojNS4+Nt*v-6ab:tuo-yEn1|CDSTWn*bCDSTq?/JwbFXfgUj56;-\\\"\\\",2):f"));
$write("%s",("(\\\"\\\"{61\\\"\\\",2):f(\\\"\\\"}=a9bwWab|5og7rLpl\\\"\\\",2):f(\\\"\\\"{<qvzWsZa7,zoW5aLc:=uVavFjT:iybn;ywP61@7VhbBWfEM.\\\"\\\",2):f(\\\"\\\"}6pKwbbtH*SszP<7Ya8I,6AbFbTazb:qebaqSOvbebqItb+bj0.VQavbQay+db*bYugb,z6;Qaxb2+V\\\"\\\",2):f(\\\"\\\"}Fah*gkRjQahb-bnyA,mF5wCg3r\\\"\\\",2):f(\\\"\\\"{t5y;67Vub;*Szub7VhbcAGhgAUqOaPt\\\"\\\",2):f(\\\"\\\"{fSqM9p6,SPqiGTaQrVP-b9s+bOaGhIP3yn=zi\\\"\\\",2):f(\\\"\\\"{wo3aAbB\\\"\\\",2):f(\\\"\\\"{Na.w>ybbub9+-b0bh?Ca,DM.OZ,bMZKZIZebGZvGp<y1/Ezoe851lbJu2bB1-|RaJ:Lu<L267CR9=a-y3O<a=uVam|xb?6hwhKwbJ3Rab;JoaGR\\\"\\\",2):f(\\\"\\\"}d.4bVa8y/9jq\\\"\\\",2):f(\\\"\\\"}bkKCfm;3bYnes4=J:LuS/PbvdOEbdRp\\\"\\\",2):f(\\\"\\\"}6JHWaW5/b.<hbpUmbOEBE<mHy7b@a2-YMJ3uv*rS9wb@NEa7C3rJ:LuTHX@Eaq\\\"\\\",2):f(\\\"\\\"{A=Oa/ps>8bl0o;GaP:*yOr@NhGY:R4R*2kp.FaJr1|lbDU;Be67CR9K.Yn46lb>:8*+ZaL46l<IuEsNv<6s7F5M4/UvbR/5MEczPhbPaqPbrQrKk1bUpW"));
$write("%s",("5/b|bl?ytJ3C=*pab7,VSf3lO<SubhbSoK0Q>|btuLB0\\\"\\\",2):f(\\\"\\\"{m-\\\"\\\",2):f(\\\"\\\"}vlC6=PfDM1H2xkbub?aRas=Rnhz.zZHTajb0b=vstAW1\\\"\\\",2):f(\\\"\\\"}I=z6abdcz91xb;su5c,sGAUYangS3uf0\\\"\\\",2):f(\\\"\\\"{xbQ<vG\\\"\\\",2):f(\\\"\\\"}vXM\\\"\\\",2):f(\\\"\\\"}vxq>arF*qWoCZHIp,Ut@JRWqkj\\\"\\\",2):f(\\\"\\\"{NJ>wj,|OlyA,?YQ7|iVGnQ<aXa+5x>Y|;1j<e1r/@P5ZQa,b,ohEqASswb;1j<9MjbcYMfqQRar-E953mP:-Aa+bN:o,T\\\"\\\",2):f(\\\"\\\"}56=u,P26TaWax6=aV5DMEaJo:uUaeb-bQuS/=vP1KAqsSjZaD5>agb\\\"\\\",2):f(\\\"\\\"}oz7?+.weEDagbMuKu\\\"\\\",2):f(\\\"\\\"}oz74s3rEU-0@a2mO*Pa2xU3I9+dfzY4d4coa2mJszo-b6b\\\"\\\",2):f(\\\"\\\"}bdV8@ijb.=utr,ls6sbQWCVq<WW.Qaab1Hdw0|a0gy;p5blb0D/F1whb+r6bybmz0/8JvfJJebgvr|?N0z.bky5bwbd+?19wAag1uoO0i5akc,|CHt0T\\\"\\\",2):f(\\\"\\\"}ZrlbWy6A+,|0:uib58x*Oy5b>aFXkuYwj,ubXamonK-,56XES0Jdhv7@/b?.gbYwkuB+LqS|RWDa*qAWEajbCgxTxquERWuZw2<nvo"));
$write("%s",("bb3bffFw2@ebIB0>l|o2>auRJ2Qiq.\\\"\\\",2):f(\\\"\\\"}i>tvb5b0bAye?lbV6>tuZw2u,h9t0Ya.Q\\\"\\\",2):f(\\\"\\\"}UNaSOjO5>G9a$dBad7cbQy8@BMAp;T>9wbpwuRJ2Zp8bGA6skdvAFXUa:>j0IsGs:9fbXoWa-0a1*q/0mbpUmbMo+b0s\\\"\\\",2):f(\\\"\\\"}GcbX*QHW3\\\"\\\",2):f(\\\"\\\"}nF-4bRwhg?UZ\\\"\\\",2):f(\\\"\\\"}.bh9V\\\"\\\",2):f(\\\"\\\"}A=.*nyW7tujb\\\"\\\",2):f(\\\"\\\"{b>t*p-bGhH=k=ZaEatb\\\"\\\",2):f(\\\"\\\"}UGKivEf>t||5N@stuoD\\\"\\\",2):f(\\\"\\\"}Gcbs>EatbUgwWmv70XrWuk=Za5bRoPael?QoBr|vDtD|bk=fbTAT-=PaEld1b3Q>adwj,UtV0Vsny0C7u>a1bN7-tq\\\"\\\",2):f(\\\"\\\"}R;\\\"\\\",2):f(\\\"\\\"}bo,Opwb91WOTa6blKgy|bhDwX>awbdbmxCH.bO9iSandmg0VAa4bpzZCVDWs,\\\"\\\",2):f(\\\"\\\"{ws*bZ\\\"\\\",2):f(\\\"\\\"{mA6<X4;sWD33nKVa.bRZVBQaVa5|Rarzm\\\"\\\",2):f(\\\"\\\"{<X\\\\\\\"\\\"),\\\\n(\\\\\\\"\\\"tb+bG;QQQr8in-<H,FaEaO.ED.UVagBGhx2lH4-ApgrVaex>Cub*z49j:Z@G;QQruH8MH2-c9U<VSZ//jH=GBEXalb|b0CE\\\"\\\",2):f(\\\"\\\"{-bi"));
$write("%s",("GtbjbJThbNE0Q2bGpSaC\\\"\\\",2):f(\\\"\\\"{R/nqRo*3\\\"\\\",2):f(\\\"\\\"}bOalbFABaH-WnScnyjbw,XM:>y1hbEQn-Rj0CP-bbuo/|@KmbX;.9RDQ|yP/M1ba0-M.-aTa?ayuFa6swb3xQADaqA+dv,h+Sazo-bhbjO>nW|e;agcvbp?WAH\\\"\\\",2):f(\\\"\\\"}WNCa*q\\\"\\\",2):f(\\\"\\\"}UgBXrlb+Bau=a<ao\\\"\\\",2):f(\\\"\\\"}:@q,SaH8zbSaLCTAqtMrT,5;5toDd*2btBI>=ua5=ufbCaAaet@X53*NdBJpJ1Irgy:Bn\\\"\\\",2):f(\\\"\\\"}UISa=a+bbP*NdB=aEa.z@Xgh>w\\\"\\\",2):f(\\\"\\\"}:ibubYa8qD7rM7+.Q7Xxq+ecbIrH8.bJy.QAa@aCwAadSAAXabw@4cjbScM.vz8I5bAqZM+bM..d<hoDPB8Tet@X@a=aZaKt=a4?w\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"{mwbco/ULn\\\"\\\",2):f(\\\"\\\"}bUalb8/5;|;5;|;zbl,pM:@Rw:@RwVFK@Oycbzbe3adaxXC8Hbe-JPQ*x5X;fbs+yNa\\\"\\\",2):f(\\\"\\\"{vf8za5*N8*1r0QoqfqwbW<h*/3f8Pt|*8buMz55NbbQZybYayb3b;\\\"\\\",2):f(\\\"\\\"{:uUaabu=\\\"\\\",2):f(\\\"\\\"{v<xCQovM\\\"\\\",2):f(\\\"\\\"}y:+NAu@.d+8wSaF7s5YqDf\\\"\\\",2):f(\\\"\\\"{v>nTs"));
$write("%s",("xbboRZNaWz|M8wSa3txb4rSwKN6:hbnX8ba;gblrCT+rcFaFoV4v=qu>yd\\\"\\\",2):f(\\\"\\\"}bcoXrd-6tXxfczz3bNS49CaqO48GaeOzFYac\\\"\\\",2):f(\\\"\\\"}M,w0<WT0f7eE<m/\\\"\\\",2):f(\\\"\\\"{F|ib@1\\\"\\\",2):f(\\\"\\\"{d\\\"\\\",2):f(\\\"\\\"}Nz2<WK-K|5bB\\\"\\\",2):f(\\\"\\\"}I9*FRt;sL\\\"\\\",2):f(\\\"\\\"{b,DaFq;Nl<xq*yxSYXML5b@a91wbh|J1jb4b<a:q4okb.X@JJ<Na2tJ32b4bVv0|7Z<a2UZ\\\"\\\",2):f(\\\"\\\"}/|9bwbAa=aurRo+ZqW|Zj\\\"\\\",2):f(\\\"\\\"{K1k-Vahbdo.*3bopDal0?yX4\\\"\\\",2):f(\\\"\\\"{b>*x-LqVvT1+y+U1QVa>1>+M9=uu5,b.8<aEaZIdAG6F1Mttbib+o>:CUeqew2JAafbF=Ooq3Na0|/bzb?NU6Dsj:;Aac,b<ajO..gjlQr/MGlplTBnj7l>?aNyeoSzApcUZtAaJyVaPaYqR*AaHC5Sib-b4Rl-:y.Ux>ML-7mPqO=h>P6b.-4bzb>/Gag7,bkTVh,CiWtbfUvbm3UOqtK9FaXaCweyq,tzAwBaRy+bST|bBU:\\\"\\\",2):f(\\\"\\\"{Ghxsvsab.>Rsl\\\"\\\",2):f(\\\"\\\"{PRUOiGs5g1Vajbtv,n5z/XO\\\"\\\",2):f(\\\"\\\"}OP6b-bdzdnRT?ab+:tL\\\"\\\",2):f(\\\"\\\"}BWn\\\""));
$write("%s",("\\\",2):f(\\\"\\\"}4bAaaTCPcbfi|Jvh,d/C<a.*/o\\\"\\\",2):f(\\\"\\\"{TXvuRbb9sGt0jHp5bbGC+Po5+kg*g+|Fa?a>@YajbmbH8kxwp\\\"\\\",2):f(\\\"\\\"{b\\\"\\\",2):f(\\\"\\\"{bAu=\\\"\\\",2):f(\\\"\\\"};\\\"\\\",2):f(\\\"\\\"}?*yN2J=QqQZagbS3YaSwhrfb\\\"\\\",2):f(\\\"\\\"{fIH6bG:x,Eaf001*48yT\\\"\\\",2):f(\\\"\\\"{*kVRtFt3UVI?2+MOubzu-yr+lW2bZawq1K2mMOYazu3b-:X|uMTh\\\"\\\",2):f(\\\"\\\"}9uUEUfUjbWakMF5@aQwBaVROa=rGyHIRa@?yusw.|8|H;fUZ.vx\\\"\\\",2):f(\\\"\\\"{w=+4b3zv4ltdbkrEz|iNsEw7bjbF5|Rkyv@+Qkb\\\"\\\",2):f(\\\"\\\"{T5Qo\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"{xS37M/bIq9\\\"\\\",2):f(\\\"\\\"}*r.ba4\\\"\\\",2):f(\\\"\\\"}pJsJr.de\\\"\\\",2):f(\\\"\\\"{QcF?9b-yCg:sQF8I-.8I2bbo*qtRqtQyqw2@06fU4z1be\\\"\\\",2):f(\\\"\\\"{L|-U3\\\"\\\",2):f(\\\"\\\"}fbT1q5PUmq9U033x72nUuo4=Ga/PGzdbT1Zznw;T*bUa<z.bjb..IgbUmo,g>nvwjb7-.boNXO/nV0Ba.>wbEaBa|bibTwebFa0t6x\\\"\\\",2):f(\\\"\\\"{|ybB-ThT2\\\"\\\",2):f(\\\"\\\"{Q-nnULnbo5b"));
$write("%s",("SpYaQq7bU*?xdbpF>afbmpfbwb8bOFbbW.VapBibnre8U4G-E-3bl,G\\\"\\\",2):f(\\\"\\\"}EDKBb4+b-4DadAO0VaV-e0xvgchK|bEwM\\\"\\\",2):f(\\\"\\\"{/glCKs6;mb=ryv;wVoBaV71MbxR?|i8I.b/qaxtDy,9b<y-bbbms+5dSdb>SlOrFlBhpcb7b0sQa?R\\\"\\\",2):f(\\\"\\\"}=CaFK=BpMWa1b5Pub1=?a*bZ6db:0d7<7:Q|faxeK,b8sC,0+Z.Y-Tp8*70NaabIp2nSIeb4bzoG->a*o\\\"\\\",2):f(\\\"\\\"{bU+\\\"\\\",2):f(\\\"\\\"}i0Czi>azo?x72\\\"\\\",2):f(\\\"\\\"}6M,Hp*b<ylbloRnil-K+OyA\\\"\\\",2):f(\\\"\\\"{91I*?2G5sOFW;U;gH6K0xM++gNaPa@ab4\\\"\\\",2):f(\\\"\\\"{bZa6sMf9bzoDQ:@\\\"\\\",2):f(\\\"\\\"{btQAvaiKOT5quOa0t1zi\\\"\\\",2):f(\\\"\\\"{J:Ca:@9wtbsGRyzzwq9Ngb*\\\"\\\",2):f(\\\"\\\"{+qtsybtqTaVsRaS3vq2\\\"\\\",2):f(\\\"\\\"}xbW3F6pQSo@aS3DAQHDaN1=\\\"\\\",2):f(\\\"\\\"}=phctvK-h9ubpQ+t|g\\\"\\\",2):f(\\\"\\\"}r\\\"\\\",2):f(\\\"\\\"{r4q=a\\\"\\\",2):f(\\\"\\\"{|Sayb,oTa\\\"\\\",2):f(\\\"\\\"}b0br@uMCwj<R:KAIsBur7Inxb6q.>c5Xa5b2*9bQ>dx0x:u@aM\\\"\\\",2):"));
$write("%s",("f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}bDaM\\\"\\\",2):f(\\\"\\\"}<s3N9tabOa0\\\"\\\",2):f(\\\"\\\"}iu|bOaabGag3i;dbGskbYNiuUaU*YNdo?6,bfbybfb?atbQr3bSD>a4bU1Thv.*O-pC.t3\\\"\\\",2):f(\\\"\\\"{tix\\\"\\\",2):f(\\\"\\\"}vM\\\"\\\",2):f(\\\"\\\"},6EP8bTa;pOFhv.bevSaS=o/iJL31w.t/bOaz7ytq?kbCz9b/b@.l?8wlbM,tby@IMe,DazogbtbosXrhJBaQr,rs<F|zPzbDa5q@3abqPlP9biu1bU1y8@nu=Gh?vRaENAaxJ+rb\\\"\\\",2):f(\\\"\\\"{Hy3bkb+y0CPa*nW;>O@|+olbJ\\\"\\\",2):f(\\\"\\\"}dbKMOaSaW5POz2qN2wuId<\\\"\\\",2):f(\\\"\\\"}b\\\"\\\",2):f(\\\"\\\"}@fbubj<-w|b\\\"\\\",2):f(\\\"\\\"}btbOa8bDa+J36roazf*hbO\\\"\\\",2):f(\\\"\\\"}iyA>zo5r5oWNs-L4U0kb9sbbV;T;|rHp86zFEar,LyEacqHpbbzuj/yb5brJTh4E0I*MAp0be1C=n\\\"\\\",2):f(\\\"\\\"}?akb8u|f@yPFNafbYM3owtj-Oa?ambq5j\\\"\\\",2):f(\\\"\\\"{Y*/jHKEa?aHC7oZa\\\"\\\",2):f(\\\"\\\"{tSN4bU+5rAauJ8bT05r>n+5k9q5wb+yhb+bgxC=@as5W|Su1HlbabQr1b9NQaq5EaDaRajb>ap6OaH,=\\\"\\\",2):f(\\\"\\\"}72.<"));
$write("%s",("tvwbs2@.lbM\\\"\\\",2):f(\\\"\\\"}vDduK-,buJ6bYq<FM\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}v2@Uaztfbh.>aPazj.<ZI8b-=57eGJ\\\"\\\",2):f(\\\"\\\"}-DFaIM=akbYa*b7zIMXtuJIdkbkb0b<u6tu-AaK|fb/bPK5MU0RaR7Pank.vW.f\\\"\\\",2):f(\\\"\\\"{qy6sP-\\\"\\\",2):f(\\\"\\\"{x-bqslvghebZs8u?*Xa?<Wn1|F5Am5G+K*q;xG8EwRvh9Za<xubdxG<7b@-db6x*r+bfHM7K69Jvx82Aw99\\\"\\\",2):f(\\\"\\\"{bQxFaxyjb6t<a,b2baqjbyb\\\"\\\",2):f(\\\"\\\"{bgb5;-t,b3b8LM=-:wbRD>1,H614LUg0t2t\\\"\\\",2):f(\\\"\\\"}bgbs-+e3bFAOy/|>a0nz*?.8i5bebN13bl\\\"\\\",2):f(\\\"\\\"}7\\\"\\\",2):f(\\\"\\\"{FKGasAmIAK6*,@5bL6;2mbw+,bVaUaI;LBXaW9xbOaPaNabwj8FANKfzS\\\"\\\",2):f(\\\"\\\"{.p4zC,VaBaVvn\\\"\\\",2):f(\\\"\\\"}jq9ubifbcb8IUIdb+bybmb+yC?Y*zoeb3bzb=aTyhbQD:qfb|J*puoB4Falqt3UahvEp4\\\"\\\",2):f(\\\"\\\"{S,D7h1*bfK4b1u6G0;.IBt9y4DUIyCM.hJbs\\\"\\\",2):f(\\\"\\\"}pM.pF,xOyQG<aPaFaib6btblI-6>aA53.,bM?Y2,xV;\\\"\\\",2):f(\\\"\\\"}bopO"));
$write("%s",("*mb5bWa,*hb;yC.PcD5VaGa:,EHhbCaS7-o+o1AAJ|b/|4bwbwouoso9+tBCxSaXaFas/Ua0rZuQaWaMokbAyv4ct=as;B|9bfHt,AuFnDnBnUay|<nh*c:Ca5n:+fcgbl3?FKrhb?aubyG<yEIQHm;jbbb>uhqhbTIzb*bpw.*Y7\\\"\\\",2):f(\\\"\\\"}IeE3*Xa1*8\\\"\\\",2):f(\\\"\\\"}1bcbe91lWaM9WaDyGx*bIzzbitgtM\\\"\\\",2):f(\\\"\\\"}Rv>xQa6|bbL/wpibVh\\\"\\\",2):f(\\\"\\\"{A+C2u3G7b>wNF2bvb13;s-b0:XaRvhsfb-b.8CyubUa.??abb|rj+tB+b6bRaX-A;W;q31.I7?aRvs<fy0wAaWaJyT05bNqVGO7FaM.whCaub?+Aw1o/odbjbAw.p>*Z0Yv79db4=H84yT;j,S*C?zbzo@\\\"\\\",2):f(\\\"\\\"}@a>\\\"\\\",2):f(\\\"\\\"}<\\\"\\\",2):f(\\\"\\\"}NG@a|b<4\\\"\\\",2):f(\\\"\\\"{<68RCUt?<l0ywBtjby-K\\\"\\\",2):f(\\\"\\\"},xq?xb=p-y*>\\\"\\\",2):f(\\\"\\\"{v3bjvu1@awp?.tbq,\\\"\\\",2):f(\\\"\\\"}n|g<nV>l5=,Q,s-Xaa84\\\"\\\",2):f(\\\"\\\"{y/M.ZE>GebhbuEj-,b.3FFOC6b*bu>+e+vPnJA8b<a@azo<a/9=aDzi\\\"\\\",2):f(\\\"\\\"{AoS+3E/;1EhbQETpNtUD8ba8;uS7cbyb.bdb7bhbgr1bawN6Ea"));
$write("%s",("VaY2k6l\\\"\\\",2):f(\\\"\\\"}ytEa\\\"\\\",2):f(\\\"\\\"},9-hbEaxboDxqwb>@2\\\"\\\",2):f(\\\"\\\"}Iov8uvMqJx5A0bk<tm=|Za2bAa3b9b+b?E+A=Ecb;EA>XaZ\\\"\\\",2):f(\\\"\\\"{.byq0rjbk96b*3-9NaXan@ab<aw6Gas*wFpsTax>N=Ya=+lyKqt^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^[2fha\\\"\\\",2):f(\\\"\\\"})3(f\\\"\\\",2):f(\\\"\\\"{#v3rga(f;)0,73-c1bTa0t\\\"\\\",2):f(\\\"\\\"}-<atbL8J>Z6.v6xXaX;FaWzywjbt<2b.|Ntl0Df8o?+lp|nWzxdTa<aQap?@a7bzbTwOtbi8nab|xjbTacA6|a5-yqz1B;ogbT\\\"\\\",2):f(\\\"\\\"{|5-h|b5C.:F5A?8b|g;tMD9bDaQqu5il1;zAy.\\\"\\\",2):f(\\\"\\\"}CQaybN:3k|glCi>yCUqutivI>JBe2ScwbiBMlK5Jq>Dnyp;db\\\"\\\",2):f(\\\"\\\"}bjb/CCa9bFahblbToQa:ogb?a0br\\\""));
$write("%s",("\\\",2):f(\\\"\\\"{cb=ambPaSa0bB7vildX3+baiq>w\\\"\\\",2):f(\\\"\\\"{mpwo6b<DQaZaZaPfnpx6=w>wvuVa:<y4m9r5\\\"\\\",2):f(\\\"\\\"{<4-MpcbxqMA>+zodbhc,-Qas++b7bHnvgpB+b?y6b+bYaYaVay4Va7b.bXupzr\\\"\\\",2):f(\\\"\\\"{Wq/bIymbbbjBhBnyU+Tak=Ra@sQaDaTB?yHpFp48PBJ:RaSaU4bbU\\\"\\\",2):f(\\\"\\\"{H<Mu-bT;Ya2b|b5b@s.bfC|0S0Ya0b4zh:W3;54bAvCa1BP@nh><RaCa?aTh+?Pz\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}xAVaMlI6SakxG8twpB/-ws>uS0?a1rbyZz+b\\\"\\\",2):f(\\\"\\\"}bIn<ambb2vbC?mw,b-tkb|-T/JB>vdb:>|bb2rz?kSaxB5;QytbAaj\\\"\\\",2):f(\\\"\\\"{BaGak3Mp;sU\\\"\\\",2):f(\\\"\\\"{/bO7;uNaRaP@Pax+?aEaZa8xIr*s5+\\\"\\\",2):f(\\\"\\\"}3i\\\"\\\",2):f(\\\"\\\"}/yfb0bwqeAg\\\"\\\",2):f(\\\"\\\"}Ir+rvbnyx/KuhBj8B7@\\\"\\\",2):f(\\\"\\\"{du/bEaI+gtB|cbEa5bMpzbn->v6bFavb=:ubSakgM4.bO79AB74brm..<a*w:7\\\"\\\",2):f(\\\"\\\"{bstzb>aOas;abFa3rS3*p?aB,pw<aRa,b3nib\\\"\\\",2):f(\\\"\\\"{b1,asjb\\\"\\\",2):f(\\\"\\\"{s"));
$write("%s",("zbibib\\\"\\\",2):f(\\\"\\\"}b+b7qiv6b3bKu/1,xSsS,|b-og|Th@0*\\\"\\\",2):f(\\\"\\\"}>0\\\"\\\",2):f(\\\"\\\"}?,,db-.r>j9U\\\"\\\",2):f(\\\"\\\"}Fadsp6Wawb+h+b/.<njyhbT1R*8bvbq\\\"\\\",2):f(\\\"\\\"}i|-bEpUaUnT.Y2UjEpj\\\"\\\",2):f(\\\"\\\"{4+QavxG\\\"\\\",2):f(\\\"\\\"{c3a3zbY2ib;9>4>qM2j/D>DpB>vbDyabcqduIrBa3vRaWae=Uja-socbmbj8X,5v..OaS7Kotb@am/F6?ay+>q+b,z?xPoibN6YjK*zbZ\\\"\\\",2):f(\\\"\\\"{-:E:.rL3qsgrUa7bG;Aa6bgb2bMsPwD\\\"\\\",2):f(\\\"\\\"}Cnk>6<q-<uCpn./b,.5bybabNp*bVae=9bBayzWa=+*\\\"\\\",2):f(\\\"\\\"{91h?0t02:xcbn9eb1-9/soZa0bEsTrTa/bZ.4b0jil\\\"\\\",2):f(\\\"\\\"{.|9/=0nTyS\\\"\\\",2):f(\\\"\\\"{*6I84t<am=X,7bI>hb,bubQ9wb/bl2T4l20b6b8r?aIydbzoabZ6-tQ*.dbbjp,/eta58bE\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"{b=rld:<jzhz|bfzab?*b;5bL+B8QaR;k8i81bm*ibRa6*btcz2kubd:UtctatYsWs\\\"\\\",2):f(\\\"\\\"{bx4Y*:rj3N:EaQoJ<OaZaS=sqdb8\\\"\\\",2):f(\\\"\\\"}ubGhj2GstbO.;\\\"\\\",2):"));
$write("%s",("f(\\\"\\\"}ibmgr1Wa5t<ngrOt-\\\"\\\",2):f(\\\"\\\"{o,\\\"\\\",2):f(\\\"\\\"}w;;DzHp+3Q=*b6by,gbX6.b\\\"\\\",2):f(\\\"\\\"}bVa-b2b7=ixe=2x,b6w7bPo1r0bUgQaLx>nkzZzq1A46bkb-=VaZzoqUaj-Bakbz9-;Pa+b\\\"\\\",2):f(\\\"\\\"{r2:30|b4+Pfp12xczgrkzUa3x@aQ7Qa1\\\"\\\",2):f(\\\"\\\"{rtub0b/lmb8xL/B|vbfiNa:xDaR*||i\\\"\\\",2):f(\\\"\\\"{WaRnCg.vib6<Ba=a.bsuAx.3wqcrziCaO4abQy9\\\"\\\",2):f(\\\"\\\"}k9Q5Xu8r/b..\\\"\\\",2):f(\\\"\\\"{bTa2w1.Qa@absubblUa-<57B+<a1r5bXrbb4bg*Cg1wngq5-bDabdhvDx7onr\\\"\\\",2):f(\\\"\\\"{babBa9bRaA5Cwc3ab3bTaDwtb-.Nt>aDw|uf8aw>qQobbkbAaBadb7\\\"\\\",2):f(\\\"\\\"{5bFao0<o,|?3ppwpnyB2,bab>aEs<m\\\"\\\",2):f(\\\"\\\"}-\\\"\\\",2):f(\\\"\\\"{-1tx-6o-wz/Mq\\\"\\\",2):f(\\\"\\\"{wS/*w24Fzzb+bIy5y1uP+?0Vhx.z9WnaqjqIzYaWal-W50/Kn-ba52bRaGyy/xbxbYaUa-ywxhbjbR6;rfgm|J3\\\"\\\",2):f(\\\"\\\"{6/bxbPalt@aG:3:Q9sy,w0b/j+:V5VaG6<68bEaR*L4,y?xN1W0rwwb7\\\"\\\",2):f(\\\"\\\"{Gae4"));
$write("%s",("hbTa36G1aqys6xR*>a-yz:Vpxb7bmb6subeb//8bXyhb/\\\"\\\",2):f(\\\"\\\"{,y8bibxb9bs3f1@|4-Xa2n?2Y8u1j:u1Eambo\\\"\\\",2):f(\\\"\\\"{Ya/ta0P/j3=am\\\"\\\",2):f(\\\"\\\"{*b7bu\\\"\\\",2):f(\\\"\\\"}Qafb6bQaSuuvgbTaKq@77bkbFztbabbbAaOrwr.rDaabIzT.V/\\\"\\\",2):f(\\\"\\\"}q:sgbCpV2Ea2bmbr+Q*@71bD5Z8NtSc-b3b\\\"\\\",2):f(\\\"\\\"{bGhyoilQzS2Box7W-5*Ea9b?4O2doY-W-cbDaYnwb57zo|bVpcbB+8bBa,b=a|i*gXaAa415bht>a:t8yx6lb,b>4G|8oGh\\\"\\\",2):f(\\\"\\\"}tW3Lucb*biwL0qwzj2/?3j\\\"\\\",2):f(\\\"\\\"{hbUa\\\"\\\",2):f(\\\"\\\"{wExjbXa@\\\"\\\",2):f(\\\"\\\"}+r\\\"\\\",2):f(\\\"\\\"}b?wEp/bw*WaE-VoN7cbeq-t0b0xcbsyat|60bh|D+B+DaR-Zty,8bT.*bK*Qa6\\\"\\\",2):f(\\\"\\\"{w\\\"\\\",2):f(\\\"\\\"{1bgh,,Dalb?au305Mtzbh1TaD5Fazbcby/mb?aNaJp+bgb0b0,U6jt0bhtQutbSatbWalb6x,bkp:sCgjbwvlb,x+nhw\\\"\\\",2):f(\\\"\\\"}qTaS0CpQupw2b@1f77bWa?aW\\\"\\\",2):f(\\\"\\\"}H\\\"\\\",2):f(\\\"\\\"}|r2bDaVhv7Brh58bH5-b/bjbub;z\\"));
$write("%s",("\"\\\",2):f(\\\"\\\"{bEa,b9bZa.b;,xtkb;29brv:vQxOaBa0b1zwbzompmp8bB,xbw\\\"\\\",2):f(\\\"\\\"{Nak\\\"\\\",2):f(\\\"\\\"}2b;\\\"\\\",2):f(\\\"\\\"{q*U+3bNaebRach3re6Dn|b2bAq2mWaTaXaR5Sa?.\\\"\\\",2):f(\\\"\\\"},WaSaVaSab6lbw6\\\"\\\",2):f(\\\"\\\"}vkb|bqwgb|bRaVaTaBqVaRa/yAqTa=a/bv,4bc,\\\"\\\",2):f(\\\"\\\"{qehp/Z.e6R*k5ZbEaSa:-?a7bu1BaR5A2Wa@aDa@amb@a2bRoPoa/-sW3,bNqAa;ptoBagqhb.drqtbx0Cve\\\"\\\",2):f(\\\"\\\"}Xac\\\"\\\",2):f(\\\"\\\"}xba5<*2se-1\\\"\\\",2):f(\\\"\\\"}KkC4\\\"\\\",2):f(\\\"\\\"{b8bUyYaa1EwGxVa0bybibOavxubW+8rgrZzVac3zbkbOazj?a4b8rRn7bmwilf5\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"}Q2AaubybQaCa.zYa+bsyEgub3b@\\\"\\\",2):f(\\\"\\\"{Oa.zM+7b\\\"\\\",2):f(\\\"\\\"}g?a3ba0<y:y?.Mt/b6ydrWaOa9bOaU|S|N2L2J2y4FndxFn:vhsF2O|-b3nj3Posz?aab+rgbMq*bwbCqAaEg@a9bQy6bhbRaq,X*dp+*hb\\\"\\\",2):f(\\\"\\\"{bR,zvpw3pUtGh|lVa?aOa*bcdSzZakbSoRa-bFa0bGvLnhbPf,bPadobbJ-r\\\"\\\",2):f"));
$write("%s",("(\\\"\\\"}p\\\"\\\",2):f(\\\"\\\"}Pi=rs0:x,yB-vbXaf1;.\\\"\\\",2):f(\\\"\\\"}wj/;-.dfbPaW-Sa\\\"\\\",2):f(\\\"\\\"{n.b@yfbzbXa7b|0q|@a>a3bppNqL|Ya9/=afbab8bYaC\\\"\\\",2):f(\\\"\\\"}Da<n/bnpmbGhTt8btbGhdtbtZs1\\\"\\\",2):f(\\\"\\\"}wb0bab;sUaCpDaL\\\"\\\",2):f(\\\"\\\"}il4uu.Q+<0T|R|AwNaWa7bfbgqhsZa4+G.|bAay/Padq@\\\"\\\",2):f(\\\"\\\"}*kMfQaFaOtB\\\"\\\",2):f(\\\"\\\"}Nalb:o+dr28bBy1/Talpfjqk/b+bPodhjbPsRajy/bZaJnybvb1b+b2b*bhbZa-bQaE-zbk|X1ebT1Na?s6w+b2\\\"\\\",2):f(\\\"\\\"}M\\\"\\\",2):f(\\\"\\\"}mv4b*0ZazbNa<vOr2\\\"\\\",2):f(\\\"\\\"},bdpgb-byb1bSaPamb\\\"\\\",2):f(\\\"\\\"},VaOa1tYaYx.reb9bVaF/D/.b60gb/+1r8bSahb;\\\"\\\",2):f(\\\"\\\"{t1Q*5b=a0jDam*qiWwk1F+s/Jn0bNakb;\\\"\\\",2):f(\\\"\\\"{Tahbgb1bdpCaS\\\"\\\",2):f(\\\"\\\"{>nqi3o4zQ-z->aablb7bIzYoG05b/bCa=awblbUaFa|b-yOa8y>aquRa4bMfHiavgwbb*gr|I*ebx\\\"\\\",2):f(\\\"\\\"{ilz\\\"\\\",2):f(\\\"\\\"}z.1uNzR+|-dx>q5++babSoZa?a-bgvIz|bboU"));
$write("%s",("aS\\\"\\\",2):f(\\\"\\\"{h|gblb>ag|vbxy\\\"\\\",2):f(\\\"\\\"}bhbrsmp@aub*gvxTqxbFs=/ebQwYaxb<\\\"\\\",2):f(\\\"\\\"{Pa0b5b0vCajhfb>apwIoB\\\"\\\",2):f(\\\"\\\"}ubMftbwbVa3b<\\\"\\\",2):f(\\\"\\\"}Qa=h9/Oa,y5/3/bo@tYahbdbF,\\\"\\\",2):f(\\\"\\\"}wmplbFsDaCavg8*cbwbtwGaN\\\"\\\",2):f(\\\"\\\"}4btbGx:tfb\\\"\\\",2):f(\\\"\\\"}bzoubZafjIz*bIsBaHiSyWaFa<\\\"\\\",2):f(\\\"\\\"}7osp*nAaebc,mbzoibSaIy2tabDaubWaSi?tDxZs/llbWaPo\\\"\\\",2):f(\\\"\\\"}b7b7b8wmbDv.bk-<o@aBaab=a3b6nltP|*b4b\\\"\\\",2):f(\\\"\\\"}b9bbt3blb8bWaVazo=a?|2b;-4e8s9oEfdo\\\"\\\",2):f(\\\"\\\"{bzbCaTafb7bDawbrucbfb1u+\\\"\\\",2):f(\\\"\\\"}ErTh|\\\"\\\",2):f(\\\"\\\"}il@rOz=op.An0vzoDaib4b.r\\\"\\\",2):f(\\\"\\\"{b5y,,xb;h*xOyybcrbwIz4bubmb.bbbwbfb<a.bwb^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f"));
$write("%s",("(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^[2fha\\\"\\\",2):f(\\\"\\\"})3(f\\\"\\\",2):f(\\\"\\\"{#v3rga(f;)0,73-c1<apz4|tbUa0b|bXawb2bBazoRnCawbGy*bAzsuMwSaWaRa@aOa.bot*bkbZr8b,bZ+TaCa3b8b-,axSaCavw/b=r.bH*cbX,l*WaWaEa9+Kslb.bEaPaebzoRa-tHt;pRa2b<\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}bH*|gibCa9+@aabcb\\\"\\\",2):f(\\\"\\\"{bPay\\\"\\\",2):f(\\\"\\\"{w\\\"\\\",2):f(\\\"\\\"{/bzoNaXsjxdczo0hebgxS\\\"\\\",2):f(\\\"\\\"{mb|bNaBnWnUn1b6rGh2o7nYwibKtp,9o4beqcb4ry+2t1bUayblbVaSp*bwp2b+bkbQa9b@aEaebzbOaCa\\\"\\\",2):f(\\\"\\\"}rIr>aKiEabb,nwp;+>acwUa1b>ambi\\\\\\\"\\\"),\\\\n(\\\\\\\"\\\"w3edoczYaAm4aO+/uGry\\\"\\\",2):f(\\\"\\\"}abmbd+,hxw+bff.bfbJoHobb0b2b3p*bXacb2b7b3n8b6bUagbQaBaEaNa|b+r>aRaubwpgyFt\\\"\\\",2):f(\\\"\\\"}nVa-rx*fb9b*b?a2blbeb\\\"\\\",2):f(\\\"\\\"}b<akbEw*yWaR*Xarw+y6b=aBvib0bRa7b6i|zOaXaVvTvUa\\\"\\\",2)"));
$write("%s",(":f(\\\"\\\"{xlbgbkbGzbb7q*s2tQy@awb?aXaOa-y=aUawbUa3t+bfbAnlxUa7|=w2bLokbmw0\\\"\\\",2):f(\\\"\\\"{Dx=rjbEw9\\\"\\\",2):f(\\\"\\\"}WafbDa5bqwktYaCaabgvBaxbEwEaGhizlbkbCsDaUaubzbZaRn1blbZzzbU\\\"\\\",2):f(\\\"\\\"}=azb?kGaVw*b2\\\"\\\",2):f(\\\"\\\"}zb<a?azoWy-bg|rkGh.\\\"\\\",2):f(\\\"\\\"}lb-bOa3b@a*rrz1wibab6bBa6b1b||wb7btbeb7bwbwb1\\\"\\\",2):f(\\\"\\\"}rkGs+bjbOa/bDa2x0b3bAoMzpxjl0u1uJmLz3yVa;hmbczO|bl3bcblbSadbFakb-y<a0bWaW|Lu=r\\\"\\\",2):f(\\\"\\\"{bfb.pBa\\\"\\\",2):f(\\\"\\\"}b=aFaj|dbbb\\\"\\\",2):f(\\\"\\\"}babCaxbXaDqbl?afb9y;pab1bhb0z4b+slb=a6b<axbMq@p1bybhrvbbbebxbkb\\\"\\\",2):f(\\\"\\\"{sgb*b2bYaNa\\\"\\\",2):f(\\\"\\\"{b6bvbQy;h-bXa|b>nrzvo\\\"\\\",2):f(\\\"\\\"}q-b9t4tFa*bnyzoG\\\"\\\",2):f(\\\"\\\"{mbtb*b+b,bOa0bgbdwZa6nZahc>a+bfjRrWz<adbtbP\\\"\\\",2):f(\\\"\\\"{Id;\\\"\\\",2):f(\\\"\\\"{4bybbbabUa5bvxFaOafz\\\"\\\",2):f(\\\"\\\"}bGtzo.bj\\\"\\\",2):f(\\\"\\\"{TanpWawqkydb"));
$write("%s",("xb4vgq>apifyPaabbtwbgb4bVnwvOazy*bmbFnkbtw=a,bSaNyYt8uFsSambdb>a\\\"\\\",2):f(\\\"\\\"{b@akb3bXaebFl*bPaOaUugfvbUaNaDf-blbPaqtNayb1utxDooxrxilsxlbtbPafjTa5b.b7bPadbvb7ztpDazzvb@ajbZa>nBa>avbRacq*b3b6b3xSawbNaczxbkx.bPabb.bNtCgwb1r4bvb<aAa\\\"\\\",2):f(\\\"\\\"{b1h.o0brvRazo+bZaDyubIsQaTa\\\"\\\",2):f(\\\"\\\"{fhb,x+w.bDaOa1bAaabXabb+rAa2b9oibwbXaRa8bablv|bWa.bXakb*bSafbZaYatbVa8bwb8lmbWa6bZa<vcyayebYxubPawbib2veydn|bnygblyjylb<rSaebPadnYo|bco3bCazo2bEsbb=aOa>aJpAaTabr3b+bcbywwwmbEaltmb?wWakb.b6b:uZa=aabib<aibdb/blxfb8b\\\"\\\",2):f(\\\"\\\"{bXazu=a1bVaXa<aJwAavx3w-bzoir-bab3wYaZaNaCaSibbCavxfbBatbgbAoqx-uEm1u3uDr@m7bXaPaUa9bQp\\\"\\\",2):f(\\\"\\\"}b9wub7bJskbmb4q.bUjGhOw\\\"\\\",2):f(\\\"\\\"{rdb5bdb0bzo*bVq=a8b;t*qEsCa\\\"\\\",2):f(\\\"\\\"}b3bYacb/bEqgbDpBaeb8bsoNa3w1w\\\"\\\",2):f(\\\"\\\"}b6bjbzo\\\"\\\",2):f(\\\"\\\"}bN"));
$write("%s",("a1bPalbAukblbxbAaxbcbLq7b8bmbCa0b*bOaYabblbib>axblbXa4e*b=aYaRabb1b<aebjb5bYaBa2bPa=rxbEa0brpbb\\\"\\\",2):f(\\\"\\\"{bto.s.bopAa9b\\\"\\\",2):f(\\\"\\\"{bQigqjbFpKkYaFa,bWayswbZaUaOautwbbbnv<qrpYaub5bZa1bFa>ukbkv=qab7b2b0bPakb/b<uvbZajbEakb+b<u5bvb*bFaebab0bXa\\\"\\\",2):f(\\\"\\\"}b/b-bZaMk?agb6b/bWaYa,b*bTaGuOa8utb\\\"\\\",2):f(\\\"\\\"{b=p6bmbBagb5b\\\"\\\",2):f(\\\"\\\"{bbbcbTa2bJsHsFs-byqwq/bUacbab\\\"\\\",2):f(\\\"\\\"}bYaQa\\\"\\\",2):f(\\\"\\\"}b+g1u.u?oBmFrCrAoEo?rbbSa*b9rXrdumbwbMt|bDa1bXa3bFaybeb5bku\\\"\\\",2):f(\\\"\\\"}sYtYaztEaXo@a5b1bZawbJd=a*bEazoUa6tzocb1b7bSi8bebXaDa0b>aSagqSaubxb:trtCacb-tbbUaYauf=a7bZaxbzj|ttbcbBa8b/bXaZa5o0bcbgbzozoSaUa|bkbzo9bvb,bRaMr.blbbbXaXa6oEpgbzb9bwpRaQalbzo\\\"\\\",2):f(\\\"\\\"{bWaBa+b3bOaAaFa1b?qQa?a\\\"\\\",2):f(\\\"\\\"{bqr4bvggb,b6bTaab4bmb0bAatbNa3b7byb@a0bwb\\\"\\\",2):f(\\\"\\\"}bzbTaFa"));
$write("%s",("7bSakbFa>aWa>qvb\\\"\\\",2):f(\\\"\\\"{r0birubfb,rXa@aas.rybydzoYaebhc3bPa,bFa/bPa-bTrQqDa.bMf7rdbFqQr7bjh@a8b|qSa\\\"\\\",2):f(\\\"\\\"{bUa?ahbbb,blb3bQaEazb7bNa/blblb+bAmVhArHmAoFmThVh@oCoXaabwbmb1bwb\\\"\\\",2):f(\\\"\\\"{b7b,bzb/bVakbNaxbppmbzb@a-bfb|b6b,bzjmb<qSaRaxbCaDa+hzbEf>aebubTa1bzj\\\"\\\",2):f(\\\"\\\"{b1bkb9b.b?aebSa2bUazo7bRaXa0bSaBaAnybbjdbcbWa0bFaSaFaAn5bOaubQa\\\"\\\",2):f(\\\"\\\"{b.bUaSaabubjbcb9bzb,ozb2b.b0beb6b\\\"\\\",2):f(\\\"\\\"{fimib9b8b\\\"\\\",2):f(\\\"\\\"}b1bdb8b.brombabfbQa|b\\\"\\\",2):f(\\\"\\\"{bUpSp>aNaFa2b@aFa+bSaEaFa=p;pvbNaub1b5b0owbPigb2n\\\"\\\",2):f(\\\"\\\"{bkbdbmb4bjbNa0hkbRavbdbCambvbVa\\\"\\\",2):f(\\\"\\\"}bebmbibTa\\\"\\\",2):f(\\\"\\\"}ptb9blb/bcbYaabPajbMohb*bBaDa\\\"\\\",2):f(\\\"\\\"{btccbVa4bZaubDa8idbVaxbDaDa3bQodbDa>a,bcbQa7iXavbvb6bcb1hjbkbPaxbNaDakb=aTayb|bSaZaFaDa1oFa.bAa0bZaDajb,b8bOaTa4b8b5"));
$write("%s",("bAmAoll>oIbKmDm/iGmWa|b,bCafbRa3b,bebYazo4bDaYadblbjbRaFa6b7b\\\"\\\",2):f(\\\"\\\"}bGaNnQa-bCaFa-b7bTaQa8nYaAnmb,bYagohofodo7b/bYagbib,bjbCaVa|bdb1bebciUaPaDa*bGhqbIn3bUa>aFaAa*hdb@a1b-beblbzb,bNa7bvbCaEahb<aCabb*bohQaub*bWaQagbSa,bEa7b6bAaEa4lrn?lXmQmOm>fXmWl?a6ghn;aemVlOmWm0lbn-bXmdmCabm6mwbic8a9mxmylRmEa0lymMl-akmIlGlVhImnlThCmAm9aAmAmkl4aol/b\\\"\\\",2):f(\\\"\\\"{f-arhubwh|e0m|mom,mwl9aEaOaqlOlzlbm5lSl6j:aqm=aAabmnmCa?lPlZl@a<a-bemim6lem8lxlamdmAa:aCa8aXl>a7l/l>l9l*lAlAaqk6l|eJlzb\\\"\\\",2):f(\\\"\\\"{l;l|l2lBaxl.l,l*bvbtb/b-aJdHdql:l1l6l4lSe|e-l3l?aAa-awl8a\\\"\\\",2):f(\\\"\\\"}l\\\"\\\",2):f(\\\"\\\"{lFa@axl\\\"\\\",2):f(\\\"\\\"{bvlHatl9a|eulxb8a+e-a1bDfqlXk8arb8a>fVhmlThil3a.iilUhQk1hsh6b-a+czbxbubHaqb6aqb\\\"\\\",2):f(\\\"\\\"{i|izi5aqbvg-aff1bzb.bfinbxbXhGh=g;g3j:k-kjj?a?e7j?j?avk2itktcBa-i|b|bvb"));
$write("%s",("6ihc6f3iEj9jBa?a-i6erhrb3bgi>jahNjLjDa?a>a-i2b3b\\\"\\\",2):f(\\\"\\\"}i;f+c/g-a6j-bxjCa3aKa\\\"\\\",2):f(\\\"\\\"{b;aigwbccIa3b1bbj,b|b0aRg3i<job:jIg-i.bPh?a=j1i/i@a-iybPc5jnhmj;hRgkjBa.i;d+cfi1a1asbubwbGh-ayjwj:a;btj1b0b-b3aAa3a7b-aGh.a:b:b,b?amhliji0i@a3arhwb+b-aPcPi/b8b1bPcxb;a;f-b0gZaNf|b.b5b-aHiti3b=fvb|b+g\\\"\\\",2):f(\\\"\\\"}iNfEf3bgf;a<b:b3b-a8b+g,bxb2b2btb;a?a\\\"\\\",2):f(\\\"\\\"{hki:h3a>a3a5anb-a\\\"\\\",2):f(\\\"\\\"{i/b3^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^[2fha\\\"\\\",2):f(\\\"\\\"})3(f\\\"\\\",2):f(\\\"\\\"{#v3rga(f;)0,73-gmb4b.bHa8byb2bhgtb=fxb5b+b<gnhRgHhPaIh,fPcsh/bHabibiFaGaFh|fld4a/aS"));
$write("%s",("h-f4a-aEfCfMaFa=alh-b;hahzhGa+bJd4h9a/b5a|fCcng-bPaBalh6aKaMa9aMaIa5axb3b.b4b0bxbzb-btbDfnhlhGaMb*g2bzb;a6e1bccJa7b?a?aobahCdYaOaVafbVaibNa=aRgRg?a;a6gVaNaUa/aRgobvbpbEa*c7bFaEa@aCa>anbJdubSczb6fMa4gyfwfuf2bsfNd3bHa?e-a/a,f:aIa+ctb,b:avbldub4bcb-biggcfgHaebdbJaGagfef8a1bxbwbtbxbUaac|b3bCffb-f-atbxc8f?a1a-a6a5bGf>azd:a,cNaGfwb.b;b>a1a,c:a-a.b\\\"\\\",2):f(\\\"\\\"{bvbxb5a1a5aCe2b-a:b1dtbHa6a/c2b3dMd-aDdBd@dmf/aob5a.d,d*d-b4b7eSc;axb+b.bbcZb0cbfJasdHa/aed+e0cGb/d,btb-b4aWbudpcgdLc=chchd6areOapc0cNb/a;bje/eGaHb5dedOb.a8aNd8aLdLa=a>aIaOaJapb6a+e5azb+cdcfbhc;aOaFdYd6aHaCa@aIaQd8aHa=a.cIbCbMd\\\"\\\",2):f(\\\"\\\"{cycvcocRapcXbocTa;b;bpbgbYdJaGbRanbQaJagbnbcb>dqc5dpbebnbOa8a0c4aJaTa5a+btb5bxbJaQa,c*cRa5a1bzc6aedMa0c3bldjd;aeded8ard5a6a5aedxb/btbvb2bxb,c1b4b3bxb1b0cocPa8aNapcMa"));
$write("%s",("gdUc3b|b+b/b2b4arcFbnc4a=a?axbtc4aSbJcPbKckcic+bZb3b-bzcXbqcFb5aMa/ancvc+b+b|byb4a9cVbNa5aRb7cFbnbFbMapb2c.aMaFb.a4a5aJaOa-a-b|b-aeb5aicybHa<b/akc>a>aXb6aOb/a8a6a/apb4a1b.b3bvb4b1b3b2b-b.bvb4anb/aJaPa5a8a4a6apbEb5a5aBb,b9a4apbpbnb8anb4aGa=a:bJacb!p@1ca61q@.ba~[2xha=s,y=z,54[54%.4[e6&yay,]99999[gnirtS wen=][c n3aea\\\"\\\",2):f(\\\"\\\"{)v]y3b&a(niam diov citats cilbup\\\"\\\",2):f(\\\"\\\"{RQ ssalc~5[~5qfa cdlnl3c/a;maertStnirP/oi/avajL tuo/metsyS/gnal/avajq5bdateg@3doa2 kcats timil.v3dga]; V);U5aC3ecaL[f6aa6hha dohtem?3e;4nga repus&3ecaRQ@3cgassalc.@6[@6ioa(=:s;0=:c=:i;)$5ajaerudecorp34[34eqa(tnirp.biL.oken\\\"\\\",2):f(\\\"\\\"{24bianoitcnufc:[83\\\"\\\",2):f(\\\"\\\"{martStup=niam^\\\"\\\",4):f(\\\"\\\"'^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\"));
$write("%s",("\"^\\\"\\\",4):f(\\\"\\\"'^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^\\\"\\\",4):f(\\\"\\\"'>3(ba7U3vJ4vba7I4.ca,4;O)?46ba5/6/#6[#6[#6[#6moa(etirw.z;)tuo.-@aba(q?b~auptuOPIZG.piz.litu.avaj wen=z|5[a7[?4:ea4302B4.BX[j47ea5283m4[x5[57gca089;/fa wohs\\\"\\\",2):f(\\\"\\\"{9[[:[[:;ba0[:[B8[j4hca36\\\"\\\",2):f(\\\"\\\"}A0batY6[>8[?4:da942>8[>8[j4gda813>8/5aR0Z0Z/512152353/2/2166263=4/3141726??:1518191:1/17[r9[?4;ca44r9[r9[j4hca21r9/da*6 T>[A8[T><ca86A8[A8[T>hca78l4.ea1312)>[B8[B8=ca29B8[B8[B8hca36\\\"\\\",2):f(\\\"\\\"{J[=8[=8[ZOkca71BU[=8[ZOhba9w5/ga141310b7[B8[B8;ca14B8[B8[B8hAU0ba^\\\"\\\",4):f(\\\"\\\"'^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^\\\"\\\",4):f(\\\"\\\"'^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\"));
$write("%s",("\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^\\\"\\\",4):f(\\\"\\\"'X6[=8[?4:#6[#6[#6[#6[#6[#6[?4~ca65&?/ma(amirpmi oic16[16[?4;*W0RB[j47ba4l<[98[98[0?@ma++]371[]591[J4[/6[<?[v3mpani;RQ omtiroglaN4[36[|U=4>[??[\\\"\\\",2):f(\\\"\\\"{UiK8/qa;t:\\\"\\\",2):f(\\\"\\\"}%%%%\\\"\\\",2):f(\\\"\\\"}fi\\\"\\\",2):f(\\\"\\\"}*-84\\\"\\\",2):f(\\\"\\\"}41ca61dA/96[j48ca8696/(a]i[\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"}+17\\\"\\\",2):f(\\\"\\\"{<84.;i:-i602\\\"\\\",2):f(\\\"\\\"{;i:911\\\"\\\",2):f(\\\"\\\"{;j:632Y:[><[?4:ca89S7[c9[9Kgca24V>/xa(tnirP.tmf\\\"\\\",2):f(\\\"\\\"{)(niam cnuf;r7[R8[?4:ca91=I0datmfB4[^\\\"\\\",4):f(\\\"\\\"'^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^\\\"\\\",4):f(\\\"\\\"'^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^\\\"\\\",4):f(\\\"\\\"'6[dM;ca38q;[|<[wHgca86>"));
$write("%s",("8/saropmi;niam egakcapn7[N8[N8;ba9tH/ga(tnirpB?[*6[*6[v3mba-?4[$6[$6[^\\\"\\\",4):f(\\\"\\\"'^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^\\\"\\\",4):f(\\\"\\\"'^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^\\\"\\\",4):f(\\\"\\\"'=mjanirp tesn|P2ca52v4.la1 etalpmet.e6[E7[NG;ba3.6/ga(ntnirbB[*6[?4;ca11yK/baf)6[)6[?4@+E0%a,s(llAetirW;)(resUtxeTtuptuO=:s c5[C6[C6[v3kdaS C&6[&6[GE<4=/ca&(?4[$6[G9[v3kba mIaD4[)6[)6[r=[&6[r=[83#iaRQ margoP9[-6[-6[P9phaD : ; RW9[-6[-6[v3mba^\\\"\\\",4):f(\\\"\\\"'^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^\\\"\\\",4):f(\\\"\\\"'^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^\\\"\\\",4):f(\\\"\\\""));
$write("%s",("'>4[#6[#6[#6[#6[#6[#6\\\"\\\",2):f(\\\"\\\"}i=[$6[$6[v3lqa. EPYT B C : ; A36[36[36[y=[#6[#6[#6[#6[?4[#63ka)*,*(ETIRWs=[.6[.6[G@nhaA B : ;,6[,6[,6[v3lba [2cF4[+6[+6[T9oia: ^\\\"\\\",4):f(\\\"\\\"'^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^\\\"\\\",4):f(\\\"\\\"'^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^\\\"\\\",4):f(\\\"\\\"' ohceI4[.6[?4[73kpastup\\\"\\\",2):f(\\\"\\\"{)(niam tniL4[164ca01?4[?43ea%%%%@4[%6[?4[%6[%6[?4[73\\\"\\\",2):f(\\\"\\\"}paparwyyon noitpo26[M45<4[<4[<4[<4[jD@hanftnirpD4[fa(f;)3D4/kaetirwf:oinu41ba2u4.ja>-)_(niamt4[Q8[<4fWP0gacnirp(C4-ia(stup.OIK4/rKajaM diov\\\"\\\",2):f(\\\"\\\"};)B3(ca11g62oatnirP)--n;n;)sn3a<a(rof\\\"\\\",2):f(\\\"\\\"{)n tni,s tsnoc gnirtS(f diov\\\"\\\",2):f(\\\"\\\"{noitacilppA:RQ ssalc"));
$write("%s",("[k4rga@(tnir>MblaM dohtem06x*3cl;abNcuadiov;oidts.dts tropmtNnra1(f\\\"\\\",2):f(\\\"\\\"{#(rtStup=niam&3kkaenil-etirwb8dva(,^\\\"\\\",4):f(\\\"\\\"'^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^\\\"\\\",4):f(\\\"\\\"'^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^\\\"\\\",4):f(\\\"\\\"'s%^\\\"\\\",4):f(\\\"\\\"'^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^\\\"\\\",4):f(\\\"\\\"'^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^\\\"\\\",4):f(\\\"\\\"'(gol.elosnoc;)^\\\"\\\",4):f(\\\"\\\"'^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^\\\"\\\",4):f(\\\"\\\"'^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\","));
$write("%s",("25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^\\\"\\\",4):f(\\\"\\\"'73g\\\"\\\",2):f(\\\"\\\"}a^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^\\\"\\\",4):f(\\\"\\\"'^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^\\\"\\\",4):f(\\\"\\\"'^^^^^^^\\\"\\\",2):f(\\\"\\\"\\\\\\\"\\\"),\\\\n(\\\\\\\"\\\"\\\"\\\",119):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^\\\"\\\",4):f(\\\"\\\"' nioj.)1+n(yarrA>-)n(=fI3c|a^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",2):f(\\\"\\\"}54,1\\\"\\\",2):f(\\\"\\\"{.^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^\\\""));
$write("%s",("\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"# qes-er()^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&/4fba^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"b8cp3dg3fw3hla1% ecalper.k4dea^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^hXc/arts(# pam(]YALPSID^\\\"\\\",4):f(\\\"\\\"'^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^\\\"\\\",4):f(\\\"\\\"'^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\""));
$write("%s",("\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^\\\"\\\",4):f(\\\"\\\"'^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\".NOISIVID ERUDECORPA3cma.RQ .DI-MARGv3g53d|bNOITACIFITNEDI^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"[tac-yzal(s[qesod(^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"))System.Console.Write($^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^"));
$write("%s",("^^^^^^^^^^^^^^^^^^^^^^^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"Put caffeine \\\"\\\",2):f(\\\"\\\"{(int)c\\\"\\\",2):f(\\\"\\\"} into the mixing bowl.^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^n^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");M3pva^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"Liquify contents ofE3oeaPour^\\\"\\\",4):f(\\\"\\\"'^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^\\\"\\\",4):f(\\\"\\\"'^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\""));
$write("%s",("\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^\\\"\\\",4):f(\\\"\\\"'3w^\\\"\\\",4):f(\\\"\\\"'^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^\\\"\\\",4):f(\\\"\\\"'^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^\\\"\\\",4):f(\\\"\\\"'4e\\\"\\\",2):f(\\\"\\\"{abaking dish.^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^n^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^nServes 164cma\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");\\\"\\\",2):f(\\\"\\\"}/****/e3a^^^^^^^^^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"),s[999999],*q=s;int main()\\\"\\\",2):f(\\\"\\\"{int n,m;for(;*"));
$write("%s",("p;)\\\"\\\",2):f(\\\"\\\"{n=(*p-5)%92+(p[1]-5)%92*87;p+=2;if(n>3999)for(m=(*p++-5)%92+6;m--;q++)*q=q[4000-n];else for(;n--;)*q++=*p++;\\\"\\\",2):f(\\\"\\\"}puts(s);return 0;\\\"\\\",2):f(\\\"\\\"}^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"))\\\"\\\",2):f(\\\"\\\"{s+=^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"00g,^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";for(m=1;m<256;m*=2)s+=^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"00g,4,:^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"+(c/m%2>0?^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):"));
$write("%s",("f(\\\"\\\"\\\\\\\"\\\"4+^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\":^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")+^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\",^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";f(s);s=^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"4,:,^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";\\\"\\\",2):f(\\\"\\\"}f(s+s);for(c:Base64.getDecoder().decode(^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\""));
$write("%s",("\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"kaAREREX/I0ALn3n5ef6l/Pz8+fnz58/BOf5/7/hEX/OZzM5mCX/OczmZzBPn5+X/OczMznBL/nM5mZzBPu++fPPOc5zngnnOZzOZgnBMGAW7A==^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"))\\\"\\\",2):f(\\\"\\\"{c=c<0?256+c:c;for(i=0;i++<3;c/=8)f(c%8);f(^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"8*+8*+,^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");\\\"\\\",2):f(\\\"\\\"}f(^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"@^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");^\\\"\\\",4):f(\\\"\\\"'|sed -e^\\\"\\\",4):f(\\\"\\\"'s/^^^^^^^^^^^^^^^^/^^^^^^^^^^^^^^^^"));
$write("%s",("^^^^^^^^^^^^^^^^/g^\\\"\\\",4):f(\\\"\\\"' -e^\\\"\\\",4):f(\\\"\\\"'s/^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"/^^^^^^^^^^^^^^^^q/g^\\\"\\\",4):f(\\\"\\\"' -e^\\\"\\\",4):f(\\\"\\\"'s/.*/print ^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&^^^^^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^^^^^^^^nquit/^\\\"\\\",4):f(\\\"\\\"'^^^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")\\\"\\\",2):f(\\\"\\\"}^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")\\\"\\\",4):f(\\\"\\\"');\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\").replace(\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",2"));
$write("%s",("5):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\",\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",185):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"));\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");\\\"\\\",2):f(\\\"\\\"}\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";FORiTO UPBtDO INTn:=ABSt[i];print(REPR(50+n%64)+c+REPR(50+n%8MOD8)+c+REPR(50+nMOD8)+b+\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"J\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"+a)OD\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans c 0\\\"\\\",9):f(\\"));
$write("%s",("\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"do\\\"\\\",2):f(\\\"\\\"{D(Integer(S:get c))\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 35 39\\\"\\\",2):f(\\\"\\\"}(<(c:++)(S:length))\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 24 149\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");end;\\\"\\\",1):f(\\\"\\\"\\\\\\\"\\\")\\\"\\\",1):f(\\\"\\\"nsys.exit 0'}\\\\\\\"\\\")\\\"\\\",0)]]></xsl:template></xsl:stylesheet>\\\":s=\\\"   \\\":For i=0To 7:s &=Chr(32-(Asc(c)>>7-i And 1)*23):Next:System.Console.Write(s &n &Chr(9)&n &\\\"  \\\"):Next:System.Console.Write(n &n &n):End Sub:End Module\")\nput=s\nprint\nqa!"));
end endmodule