module QR;initial begin $write("%s",("Module QR:Sub Main():Dim s,n,i,c As Object:n=Chr(10):For Each c in\"<?xml version='1.0'?><?xml-stylesheet type='text/xsl'href='QR.xslt'?><xsl:stylesheet version='1.0' xmlns:xsl='http://www.w3.org/1999/XSL/Transform'><xsl:output method='text'/><xsl:template match='/'><![CDATA[write,format=\"\"%s%s%s%s\"\",\"& VbLf &\"(\"\"\\\\write{-}{txt}{(\\\"\"with Ada.Text_Io;procedure qr is begin Ada.Text_Io.Put_Line(\\\\\\\\\\\"\"print\\\\\\\\\\\"\"\\\\\\\\\\\"\"STRINGz:=REPR226+REPR153,a:=z+REPR166,b:=a+\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"2\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"+z+REPR160,c:=b+\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"8\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"+z+REPR165,t:=\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"write('implement main()=print(\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"BEGIN\\\\{s=(\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"d=(\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"(a#include<stdio.h>!nint main()\\\\{puts(!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"&3dlaiostream>!!n(3f5astd::cout<<(!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"class Program\\\\{public static void M93a@aSystem.Console.Write(!!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"let f(c :Int):Latin1=if c=127then!![2aba!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"g3craelse(string_of c@x3cma g caffeine s3cba@,3oea!!!!!!!!Z3dra)@f(c+1)in print(x3ctaQuine Relay Coffee.<3dmanIngredientsu3eja!!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"@f 10r4igaMethod*3i%a);let g(String ->[])!!!!!!!!n[c;t]->74idaPut05wpa(int_of_char c)k6euainto the mixing bowl44klag t!!!!!!!!n|_ #4ktaLiquify contents ofQ3qeaPour)3w54elabaking dishL6fiaServes 1H4jeain g94dea)))sk3b[2cca!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\" [2bw3kparts(nltnirp(])]~3kja.NUR POTSx3k,3l!$3zba!!&4l!$3lJ4nda[))r3kq3mL3k!$3|[2\\\\{ca\\\\};F3Aka)1(f\\\\{#qp]\\\\}Q3Dfa3(f\\\\{#K3Bga7(f\\\\{#.L3Bca51>4Fba105Gga36(f\\\\{#\\\\}6Bra21(f\\\\{# D ; EYB RCb;|X3(da,43O3HdaDNEE4[O39da. A36[O3<eaPOTSF4[46=36[O3:maRQ margorp d6HeP4[O31baS;6[O3;A4[JC2ca52A4[A4<ba&m8[C49gaS POOLoA[O3<ea\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'&,)F4[oA;ga. TNUO76[O3:fa(rahcr:[96<gaB OD 0rA[O3;ca&,C4[H=8ca)A|8[3?<eaTXENz8[z8=66[dJ=haROF PUDK4[jJ[%X[K3hla(f\\\\{#(tnirP;jZBca76M;Owa;TIUQ;)s(maertSesolC;)W4C\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'8Jla115(f\\\\{#n\\\\})2i3aL4[683da201C4[O37ia402(f\\\\{#\\\\}D4[y:3ka904(f\\\\{#mife<Dh:Kda918i:cj3bM4[:63ca443@[86:qa811(f\\\\{"));
$write("%s",("#;)\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'\\\\})8868zCGT4Mfa30603F4[@69da526YVaja,\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'&\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'(rt.\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'n<[wC4ca14&8[g<:ha722(f\\\\{#pL[;53ca83#8agaq\\\\})677q<a;6[\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'86ba6C?F:6T!$8[qC4ca29s8[qC:ia07(f\\\\{#\\\\}\\\\}6H[w8[D4[D4qyTaw8[3F7ba9&?bba4:6c96[bW3hL[Q;;ca39QBaj:[O;;ea&dne>=[O35ba9)F[R39da954MKaz8[z84ca9506[*?;ba4)?[)?Cca6396[*?;ba7rQ[)?A\\\\}a&&PUEVIGESAELPn&&&&1,TUODAERs3ak5[XM3ca80;8[YM;ca45;8[NVBea0658:6[F5:ca87F?[5Q[D4[PFrca705Q[:5:ca03:=a%a&&&(etirw;\\\\};u=:c;))652%%)u-c((||N6[88[D4[D4nda43388[E4:ba0PHaEJ[iE>ba1hE[hE;ca73kPak:[D44ba0PQ[w8<k:aga&&&#-<46[*?[D4[?=oba5Q3az8[F46ca83*?[n:Cba2+?[A=<ca16k:[qWBda||imJ[465ba6.QFvAPca78\\\\{8[PVBea6335:6[%89da501+?[LD[D4[i:sda582t8[t89ca35lJehaBUS1,OD96[#8[D4[O3n~8[R3:da990.?eda944+H[v::ca98.?"));
$write("%s",("[j:[D4[lZu|Q[mZ=ba4.?bta(etirw;)3/4%%i(&&&&i4B/8[D4[-H-ca39.8[v:9da307KV[F5Bba2N4a96[R35ba6!$8ai:[JV>gaESAELPL4[??3ca44|8[rC:ba9pSa\\\\}8[LV@ba1tL[~A;ba2hLG:6Kda991qAG/6Nba7KMaj:[,?>|JbQa\\\\}2=:/t;2%%t+2*u=:u\\\\{od7 ot0 yreve;i-=:u;1=:+i\\\\{od))1(evom(dro=:t elihw?s;)s*||B5[3Y3ba03Yar9[#@5da533s9[~@Cda960;6[@W;ca65~@[pR[D4[-Gsca28s8[ZJ:ca18~@bha#-<1,OD76[\\\\}8[D4[+?oJ;G\\\\}8Oca37\\\\}?a3W[O3?gCa:6[LL5ba59Fbk:[gKEIMC*PKca57~8[95:ca65~8[LD9ba8>UGMDP/6a.?[IU?ba4Q3a:6[\\\\}Y6ba8~Q[.?Cmbn&&&&dohtem dne.n&&&&nrutern&&&&V);gnirtS/gnal/avajL(nltnirp/maertStnirP/oi/avaj lautrivekovnin&&&&R5[~R3ca19&9[I>9da917&9[EWCda586:6[nM:ba5%8F&R[D4[h:,da734s8[s89ca10<5aba&[2aeb\\\\}\\\\}\\\\}\\\\};0=q;)]q[c=z(tnirp.tuo.metsyS;)0(tArahc.y+z=]++n[c;y:]q[c?n<q=y\\\\{)0>2%%++i(fi;48%%)31-)i:3c&as(+87"));
$write("%s",("*q=q\\\\{);43622<i;(rof;n)rahc(+g8[L9[D4[D4otP[R3:ba0tPbgaq\\\\})299:N[7D<.Wa!$8[j:[D4[q?oba5tP[CB<tPaW@b[2c=6[\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'8[D4[\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'8oba9tO[&8;ca46wY[#8Cba5nC[nC;ca88i:[vYB[2goa=]n[c);621<n++:Jaqa0=q,0=n,0=i tni;\\\\{5[\\\\{E3ba6JO[)Z;ca61U?[?XCea0632;6[F5:ba0.LG\\\\{E[y[=\\\\}7[R38mFaT?[Jc&6a2b9aV.2a4a5azbud;axbs.54k*Ga6a2b5a?fLa4a/c@cPtK6JaJa?f-acVxbwfzc6a/a6aHb<b<bHa6a6a>a9a@a3a?a7a|bKaKa95:aV+2aBtub8aucVjm./apd\\\\}fLt5amdfbFhpb?abdZcXcVc1bTcpcQc>a>aArzz\\\\{f3b+b\\\\{f+b9bPa\\\\{f+b8bLaJaKa8baL>a:aJaJa8bTacXJaJa:b:aLaJaHaJaJaLaJa8bZBzz3b\\\\}bu3atay-y-Ta4bzz;ay-Ta\\\\{f+b4boazz9bLaMa\\\\}bJaNaK3qea\\\\{f+b>4ae3aY3cfa8bzzwl4d1aJaQaE>;ay-Ua:aUa:aY\\\\{/apd8bMb1btb-aXcvb-a1bTc:6acawbh6a)aAr1e6a?a9a>a3a6a\\\\}bet5aKaKaBtucVj*b*b>6cla8aubJavupbC>6bCa\\\\}bUcScucVj/a.s6aE"));
$write("%s",("a9aucHh/a.sub8aub5a/bxb1bJawbpcQcHa6a/a.s3b5aJ4imaUcSc6aub8aQc|4aU7a4a<bRckf1dHa?f;a/aIduc?u8aQc/aIdHb|c8azc6azb9a2b9w3beaSdQck3cka/apdxbvbF484acaHa13gbaS/3ddaSdS/3n;apbocxdvdW\\\\}nbJazbHa6a-e9a-e7a|b9a6aQc<b=a-aztVcNe1b6a6ao3ada|b9i3fDard7apbTI,d*d|dzd5amdBrtfBe+bNrcc7aTI5a2bFhMaztVcjevbJa>a2a:boc?u3bkaxbDbyb4c6a33kKaxb1bF4vb4c/aId=a=aSdQ*Oa-aQ*OakbX5Xa7r5dFd7rDr?a4f6r4a0eDrAh@f|b4b0b0ey3cea-gJe#5azbreAi-b?iceDuMrCw.Bs.2b/cPa;aBeld8bfbpbfeubFcWbfv,bnbfeyeicefyejeJ24f6rlmEa?aMsAl<hKo>a9a7b2cye8z,b-bKo=a9a7bubxbs3e53gbaA53lG3a53gjaZo<r9a7b+)3flaNwAaY-9a7bw-3bmaV\\\\{XbM\\\\{>i-bKoi3auayexdvdtd-b3p:f-bMm1rd6eraOitrtrtr@h=j/r,r1<6diaqo-r*r2ru3araJe0e=art@h1b4bNe1L6fgaZo/r,r13e;3giaDr9dqg8e%3si3yib1rDrJele:b2f@fZ:V.2a2a5VBlog?fFrgftf0eDrp98aDrpb2fErEf@hJarcJa7bBlH"));
$write("%s",("hyeZcfeBlogybhhBl<rJaDr7bAh@E3d=3eua9a9b9a@aCaBlogyeDr>as3cba@s3d-ap9:a|b9a0b9ap97aDrp9Ia|b4e:a9bJa0bBlogXsW3c)a@aCa9aCaAaJa9bBlognbcf|c6areVjBl<r0eq5g1a4eMttbye>anbfe9apbfezttsloye5V*b.bbbye5Vye7bq3ema5VnbfeAh@flc(>aca6a,4a8a8b9a7b4eMaJaybZsg9>aJaVcrgpuTc0e<breIecf|c,bA\\\\{>aJa-PI[R39dab-ae5c1aDrDrp9<a2b4e+b|bxbvb:a>a>arc4e+b*eJ2,b4b-b\\\\{cN:ecaqn*:3i39ca4rr@mc=a(4[i3[U=%ga;A\\\\}ePmn4[i3[=5)5Ebbahn4[i3[i3[i3[X:V4aawbtfDr5VI\\\\}MZxd5bxb=ururgpu@uXras=u\\\\{u0tAu0uHuusw3a;cCsJVVvJVjXhXNU@Wgv?y5Rj+U\\\\}@WaV+\\\\{lR@WSvRW*O.9sv5VZ:lTNWLWEaVvHWzX=aT5tLHw@WuV5D\\\\{wQ*8Wp=Da8YX<d*A,UNO*0bM7wb1bYHX9Wa=aSav=zwf:,bcEnL|Yzz*bp:+DCa1EiKUBv6jbd*h1x.|*n1Va@aibv=jbXwE,h@5.V<h15D2vbypUmbZTybzbn\\\\}6+Ta\\\\{w<a?aYajbvbkbqM*bPTV@q3a7e06Ya-bL,|5|yHv2bTa:TVaEvmb>Ve6kvhckVe6kv9blbdV;dWU,"));
$write("%s",("b|506c\\\\{\\\\{z\\\\}b>Vj?J-H-:?VH9vRawv=;IvP*-b|5Jy:6SaV\\\\{bvjbI\\\\}MZ8U,?5U2bUa:UCa6H,Y\\\\{UVv;|,Y6+n\\\\}hcRupUxb|YzzpKbbGvMz;zbblbmwdbWTjbZaax?3PTV@LTpvnv0\\\\{Avn1nv.bBa,NP\\\\{db5DNa?3z<dbNvYaCa3b@at=hbT-dbEaT5tLcz5RNU,?nv\\\\{bAFXRwv4w?>O|\\\\{wywPCWaC5hb:|*L|.l-bxUu+S9553=a+v8w>:hbQdhO?>C\\\\}HwC\\\\}sY+vtdC55vxIPuEO=ajbsY+v+b7w9\\\\}+vUy:R95-,2,cv=ap:hbhb3yQ5dxM9I\\\\}MZx1CRhbY-?yDwPCK86M1273a\\\\{awzx.uApE*L?Sbwlb@Haw1,YVY\\\\{p4aGa=<URcz:/9xwRIYc9uT2BxxvxEz-TGQq\\\\{iy?QRak=CzjR?QRaYvNvJCjDwRp\\\\{:?nYr|53eGaE9jJ2Blb4@\\\\}05.4yKVRafS/S5I<\\\\{vx41zQDQHzEZI\\\\}MZm\\\\{zQI-\\\\{7-Fa1yy=O/bt\\\\{-H+3cuaPCC,A,R?f.jyT12B:40Ec3Q!$bEwWwyb7bvFv/twvb=a35,zUJf3XJI4/KhbIVX<3bnzhbVavFcG\\\\{vab95,6<af|Zx4\\\\{<af|hbK?KV7we3eb|Embf+C*35fz>a9xt4I\\\\}MZv/zOmbixt<Aa@w\\\\}5U7a0EZX/b33:Tbygb|v/:/Sz.7bL;gbCxRTm"));
$write("%s",("baxfRXaz.7bR/>5fN/3[/3oeaI\\\\}MZ33\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'Zb-X<M>Z3Yf:4;.|lUu6dWu6GU\\\\{*>aU+?SH-T0hFC0Qj|Ea,nLQ92zISnwP\\\\{kwVDeD\\\\{.IvT0hFtbcv*O4bq:qz*.v-eb4bq:e|Daz85QvEGG./DEtwmb5DGalRKEkEuG.Q\\\\{.Iv-GlRb6-wNxq;.N\\\\{MM,I\\\\}MZ2B66u3Z\\\\{NUbBrDfRGx2>aac.wEE2w:8LS.|vdsTpTKuxV,vU+3-e6:,bB\\\\}XjWi@m1Y8g6X>tHzbVbHzEZAQAZiR7bP\\\\{fbG.DYG:.VDYGZ4Q5P4QZ4CAk|:1lUt?I\\\\}MZs\\\\{6z\\\\{5fRV-q8:JcbJzR\\\\{y\\\\{Rz@Z;3sZI3z0AaRw>@KC6bHIrDCI?Sm1j+M?dbTajRoPZ2fR53a+gsTXQQPZZ?Swbzb.Zs.z0m.:1VxEJCYsOo6*E;TCv7/8PbbebabCwpM?a<TW1SBUZ?S7NK.9V5VZ:a5TGv7DYGZ\\\\}>k|.Nv:ZaRC1,8788uG@S/9|v33xv|*b6-wC=c\\\\{Wa2Z@Sww+b\\\\{.g0XaX<ixX81,/|0\\\\}\\\\{bTaQGK?Va4+*LW|5ZuybB\\\\}XqN=|M,,xp\\\\{oWlRL*JDJ\\\\{VHJHXum9iK<*/RP/wbqOv0c\\\\}v0c\\\\}JzRaP*L;08.,,,m9-X<MsZ99,XEa8bZec9lb?aI\\\\}MZX01|Mt8.2br\\\\}<wP8a0S0|R>vUai\\\\}0ENUK<>"));
$write("%s",("@ix,:p||UJ1jUexF.CxzYL.cXmwVyOdQatb2br\\\\}4bdbd\\\\}J;PTR1B;bx;02*<MsZ5>W1SBtMpB:8LSr7EZ14@QETv0u9n9ZaXab.EaAADZhRvWeI?/lV4OI9@xTaDxQwb/1T5VZ:iP\\\\{2y2K1X5Was\\\\}K;f4ebo6yR\\\\{bTa\\\\{w;WIZ\\\\}1i@VxWStVP*3+H:oQU\\\\}bB\\\\}Xt1lbpw1x-b9YbBrD0w/bxVO2L>\\\\{buGzbbB\\\\}Xz6x52bUL>*r\\\\}3:jMSB>6yvQGRZG.);acawbE;aka\\\\}9?KI\\\\}MZT=)9a6b\\\\}>@aj4*E57SBORSaT-S9V6FESV.b|3tFFa*bVaSx46c:n*G1@aj4Ua4?P\\\\{yb<aUamx@/F.\\\\{bKXZau6YyP6-A=w0Lyyv7-vrz=a7+X*j-Ua6:74Qar=eb>a3TH*y34|mb\\\\{:QaVwPaR4ajam1G.g@PB<-=hGaYZ7bHI=CI\\\\}MZGvbH?S|*i5rvSBsCF:le4bc;m1E9jJsCHI=C*M5bK?>vevIW*bL4Q\\\\}/=a?a-bO4:4:JwbY-.B+b>:.Qw8UF.80y3S:?1vo81X1-,=HwW|5Z>v+NT4m1Y8*6aNa0.9KvbavYHJw97*bkbbbybzbo0VxI\\\\}MZH,T+SBsC0zFa3btW-F<a3zOXFzfJjb4YvbTa1JNa!![2iba!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"o3j[2|pa\\\\})3(f\\\\{#(tnirP;)R3Fqak\\\\}SBsC/bm:F>QwNPo3aqaDIBJmEQPmEBJmEE\\\\{u3a|b<Z|TL;X-PODau6\\\\{b7bP\\\\{txhxBJmE4bc;hFBaNa*bb6mE5QDv6bm|8z0b1JDaI\\\\}MZUaDv.b:?,bbxvEHDVx.TkWKG=aAFVx.TSH<vLwJHDXHHx:KwIw)7afbxw,bbyL?>:zbbBrD2x1X?Ct\\\\{\\\\}/DYGZV\\\\{lC9/7bOSO|fRAaf|2by3QaeD5,k-ZAlRb6tY+dc<c4g@ZAm@PB88Ta*EwbJ?kMaeauQ\\\\{bcCe#a/9|.:9\\\\{yiZMtHw3b7vcs,bWzOZ+DBz\\\\}Ca!$bJWvb0LU6rRS;-bLSl<ibO|Yawb\\\\{b?\\\\}\\\\}\\\\{K5G0\\\\{+8U>vlbUC,OV8ZwIG9TK5b/\\\\{Z2xxPEVn..b/6+GYa4b7Kp18r:9P:wV3zXHbb4b?yp1O40=YIs7i\\\\}wbUaF4a)cP:eb3bmKI\\\\}MZ*b<aAFfJTai\\\\}bDr|+bv7-bJvi\\\\}a1RH3z,blbu61xUaROzP3\\\\}9Lj=kVe6:?>,Zwix0=YI.bZ2l-m+-\\\\}0v.*by5>T9wbUa.L-bz6K?\\\\{3vbp:\\\\{>P\\\\{87vb1Wnx-?MwE|0yp=nxu@MwlYLwsG?Cez\\\\}J;6+<|Th|T"));
$write("%s",("1lO\\\\{yyR+byQ@/5.D.Y,P:4biNE+,OC/AFG*cv4yr;dbT6cQaiDJZbRRz5VZ:UPtM4Zo6hS78cbrP:|FQO|GBuHjFZ2fRAaOyn*v77bzbTaF84-r;ext102SUOaV,cGama?S1bhb-biI\\\\{bk3a/au62b\\\\{bUVPGXaGalR\\\\{bY\\\\{*b<aWX7bhb?v|Ta?X-;VT-L4a1aeb1xR|u@gYG;jZebWaSSzbmbM?yveb0GBA+bJuNaO|Yat4acadOt4cCcUaZIEvaEC=\\\\{bUVcUI\\\\}MZm||byv.LbXS;@Lj8;Mj4mXVatbowbGU6T-5FR|xb+b+?V*vEGxfbz4iI/bT-8z.|xb+b,bb\"\"),\"& VbLf &\"(\"\"bcb+bJu2babdT.b54bb0vSX|UZ>cU0y-UYafR\\\\{b0bFaxbp6QEezYayb\\\\{bY\\\\{n*v7cH|-5:L6+bpw\\\\{5<x>?P6ldTaZIG1L=2IXw1ZEct8\\\\{bf+z4xVM@oVO|YaJDT-8z:1E<bX\\\\{bIMt:gW>Ly\\\\}xb13adbMvkb\\\\{,v/ZAlRI\\\\}MZ.bN/-U.|b/Lxh8e6Mw7bVbZacb/,c7PygzevQam.I16bOao81X;wK@9B+WUwtYa*4ZSa.bPaqEs;cMaY9NY;??U6NUaJQS\\\\}a+|TuMf\\\\}UajU/bI1r,,X@60N*b.bGDHIrDx\\\\}DI8+CJW|5Z.Bj*Faxbs3i3c/cLXfRHI=CgR|TI\\\\}MZQ+8z.|m1;S8z.|wbm*fRf-0?xvH177"));
$write("%s",("TT?>R?NUlbf:/P=CgR2bvb,b2-4QUE@LG1dB=.s|bbib\\\\}>wbUwrvcP9P4?c>3b@8QaSaWaZIP6X:;=<\\\\{,XpDH>mBH>6>b.A+WSRGb<I\\\\}MZ0;rDfRHIrDvR/bWzOZr+3P3BESSXvM37ASc4hRHEs\\\\}J5SPhDGZ\\\\}>wblbk70NTZrO?3a=a-Fo63>;WIZ0wW19VsNx|\\\\{JyQDa@8VxEJ5VZ:9+VS+0oWlR@xQY1E981WI3auahcbQWa,bWQ?Sm1-TiXTz+Ia2bHI\\\\}XRONa.Zg@PB88KQKu,eNSZI7Co,wR8b5+9BLBn+0xnM5,Ta,C\\\\}15+8Wb.@6I\\\\}MZY-9PLB,:C=6B@80vSXvMkCQaSah|zBZAsBiCcNWRYHFR2>YUk0?a/brRoN/CmJY>H>>Jaoav0A+.Th|C-O4r9r4aSa3>;WAQjRtT\\\\{Djv,?NGI\\\\}MZExO;c\\\\}WRWaPaWaO4iC.QYa,QDD8bHI=CmRz+5,Qa/brRdRMz:W5,m.dWUQamaQPmEwb@albvE|4coay-Aa.A:JAa3b5,L4a\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'a|@LzNBtbZ\\\\{1|2bmJcC+,Qaab5,RaWaAaZBl:a,byy4QI\\\\}MZX+TZ2|c>WaAa0.lvrK5D2viFQ9LzTEmbY<;2.b>v@xwxCD<M,AOaAa\\\\{JP\\\\{bbnRvTuZV9H@Y9NYzbVQ7b<V|7axL?4Q,EWaCIUx<v9JG.vdsTKZEZ1W,7ub+9aoa,b4B21I\\\\}M"));
$write("%s",("ZQzwvoGeeak-n333c9aIZf..TmJF>i54OI9nRa6*b4QESSX2Ig\\\\}iXi*465X,vU+,@-TWyTa\\\\}7acb|/.Tk3a2M,2BPy0=9FV9BB,zdT9bq:zYI\\\\}MZDaMvlVrvSBUZ4Zo6HUixczi?RaWaWa3wtySaAaOaA4Aaq9Va-c;4N)MAka721(f\\\\{#,43zNBya201(f\\\\{#(ntnirpn\\\\})215(f\\\\{##OBT4S5bPWaWaQa2=ZIp:6CF0w|z|Ua<=aLz;4O?QA@ParOeb<FZI5ZjNf:E<f|mbm*ebvU:?TCCamBQ7GaiYbB\\\\}Xgb6bmb=I6by+5ZX9Wah|+bEBUa@aHI\\\\}XqNG.QUFzp=:?-,svI\\\\}MZJ.&8e6b;=o78z9CcEf?Dv?Flewef|rzd\\\\{b/\\\\{Ze|VaYa:6Va1b,TJ\\\\{0R7bXa0=9F79ADm.F,,bxvyyO|H.R\\\\}.AO|Dv?FNU\\\\{bN+DOe:Xw337bXaM:RaFVT6Qj00|\\\\}w57bryL?>:|TW7X-zT*b+5eyaY-leQaSaPVJVVa0=cE>L4ZuR@Ra(dn*4@FLH3GQg>|8\\\\}va\\\\}UN3:KwwbjETa7bOaZOQy6zxdSYRaAa\\\\{J@P5DzvEatw0bf-3JYa*vDE@60NYZ,ZWKnv/wBF7I?vh,cQc\\\\{Aaozkb7+l:|FVbrRS;u\\\\}.0K;R?r|avXLOaN*/.?a>x6,5.KR>?1bc7O4YaybzbP\\\\{cbM@eIwbUaYa+bp6Za9b<vr9O4>zGxz6"));
$write("%s",("Dau6ybzb;UvbbV|@Lz/S6FRzPap=I\\\\}MZ4\\\\{o\\\\}0=cEsHNUV<4X|v,QSy.>MxOYe:O4vv5\\\\{/yxvowbGibx*6blbI\\\\{.QN+wKcv-Q|4IWxxmIasa.bz<cbB>QG\\\\};zz*bI1WYafb.Q+v,Z,ZxO8.BF7ISSZXlY2IezE5I;8z:DPYu\\\\}HIrDfRWO6M1bBAO|Ya2bA,nW|7M?@xc\\\\{3bv7we12ebBIdROy=6oz7bUKanbz<cvub8UpEPapM?ar9O|:T|7M?2\\\\}Pa1bLXZIP66CdM7::?-UYamViFc+|716CanW+b9.6b\\\\{br\\\\}vwF,jbR?\\\\{w;W1W>:zbc4g@r\\\\}/vRVa[aK@W;7bs||bVas|C*9.C*T0p\\\\{n<4zWzOZpF-vmF334B21>ER\\\\}i:33r|4vhVO|CI?SI\\\\}MZwbyJWKnvO2>vm*9Y5RKKaAcp:3YtbF2<aMz\\\\{bbV>GYU?aYJexEY>B3<+N7FHWm:.QMv44jSbD.vT7x|Ey4v:T2bjb2I/0Da+:B;byuv4QF>Y-Ey\\\\{dX<C,8|t|S4SX2IDaT1ASwb1bQ*iFR:GZs|3bD1F2lbubSa=aAaUa*\\\\{.bN4CaAa*Bsyfb\\\\{b6bOy5bezjXezI\\\\}MZfbBa*:qzC+uSzbOyv<NdK*Va4Xxd@|Vw5++bs|?at|T2\\\\{dC3KuRaxb/bw>O3gwayJ,Z,ZR1ubn+\\\\{dcbQRjJASa5aea,<|.IQacabMXABla(f\\\\{#(tnirP;E"));
$write("%s",("CB;b3(f\\\\{#wb;65bezNT+bdx,Z,Zlbwb;68zOy@a|.Ta>?ubSaXCG1BKI4R;ABmKCa6,E@OVYal-LVh:yP>PI|L?4@0vSX2IkC.Q@Lq+yG2/hZI\\\\}MZg.,bZ\\\\{C;,?H.ZaSx8b54U\\\\}+N7Fyb\\\\{bVDi9c!$b36=Fzb>aF?0Fle*5\\\\}KNRE5xKT+SB2By+5ZNUR;le2>YUmJ3*0b\\\\{w6.v/R|lb\\\\{bKQWO,Z,ZL?K.SB>6B\\\\{h,cQE,h@5.3bK5|TuMwAB;bylXZaybI\\\\}MZb6fHg5aGa37ETbD.vd>0=cE0*fN4v9B+NT4fbXyXa|bxx,X8SfY3<;wN<<\\\\{,X>SEJAG>xO|W;W\\\\}C=acar\\\\}S3czbAS2*<M>Z-,G>I\\\\}MZzb+Nj>SBsCnRa6GWX@?>O|W;+b>:zbbBrDQvHI\\\\}XjWV-\\\\}Mwy0Ft44xY|VQvbYx;87bs|CalzQaubG.w3?a@|-LNUW\\\\}fRa\\\\{pJD6at8abdcGR|C7.|h,a@gRw3-blembgT0vSXdO37lO?|m*i.MtcXlbtb3\\\\}UNr+I\\\\}MZ<K|6T12BlbP6z+bX\\\\{fP6z+?ayO;dbb7|59xb2\\\\}>vD.X+p|0=9FW6=27TW7cbbD.v=a-7+7+bq4f-Q0hbUabb<w\\\\{;59,b;dE5C,KY;6E>,x6\\\\}a:,b;dbbH902JwHw0B>vJz.v.02;EabXwb3b?>t4Q\\\\}IwDYG:?aOT+w\\\\}Z,Z,ZXRdTP*4=m1-T4?T"));
$write("%s",("-90lQ|T+05VZ:HFETgZUwFTagc\\\\{buG-z+zC7y?B>pxSX@|DaX-Z6lb4\\\\}IR<a98IZ<?VatbowOaZAlRm*ZIP6aEn+f8dG:J>am+n+z>ku.A84JRRVj-k,:JVx.T?K3bW1SBUZ/bxVv:Zacbn;9BGxf.WS9|hbmbk097/BlR5MI\\\\}MZxz1Vowk\\\\}SBASLX>SEJCY\\\\}Ke*c*lVrvcP@ZNRcgaA+EJbRoSaebKZEZ14@QsC04hRj>9VsNGx7Tl8SPhDpZSx@|P\\\\{87<S.NKujWO|1AI\\\\}MZA<V9wRvbRa6S4ZYZ7bSa?>tvN9wyA\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'tnirp*P[4@2ya8361(f\\\\{# wohsn\\\\})2575(f\\\\{#0B[R35da442E4E>6Tka;)\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'\\\\})00611<6[R39ea0603F4[R38.b93332(f\\\\{#\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\',\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'&\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'(rt.\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'+EJCYUaGBuH;wt\\\\{pBPu4QzTNa;\\\\}Uwd,wvC*m?|7>@sG;@3bN7|y3y:8LS.|:8jQkbD:Mv\\\\{K|8+bcEE,FR0b7bXa4HBaNaS;ub6vb.|-5\\\\}bwib13aea\\\\}8k,/3ceaf0+G+3ageg8eYVa4\\\\}0bf0b/1T,AR2iIB>GBI\\\\}MZN@V9v4TGgE5:=Fxvfb-1R\\\\{s\\\\}*L84<5b.|-N/t:gW;w,=S0|vk,s/"));
$write("%s",("mVg<OwK*v8k0WDFM+b0bWZBaO684=FuRUaiL4ZuRUa6ZrDCI?Sjb;W1WTz4bZ3hFTaAZiRSPuyL,3P3BZ4CA5bRZO|i\\\\}71NUVQXHx\\\\}8rl:nJi.|yLw957TI\\\\}MZjb;::?OeNF>EiNUD2x1X>L?vlbixczVQFc267|\\\\{@tb2xY-leX\\\\},bcXmw:9ox0=cE;w:3Nas.;UdR/\\\\{h\\\\}U*v*6blb:?csYar9bD:9tv@0NY>GWXCvN\\\\{lzjUlbBarKG.yyP\\\\{<wtY-RjVW\\\\}:T5RyR3br7QBasa>6A.H0y\\\\{Rz@Z;3sZGhy3eze7bI0=1I\\\\}MZt\\\\{PB88.Y5Ds4UNPueY,?T2mIb/DKl:<aVaQaYtrRHROs,6vbMzR1B;by@vX+z8Pa5/Oy-c>Pc<lb4\\\\{LX0=9FCBr\\\\}TChxmbB>+ePyx\\\\}V<T2f-l-.b\\\\{.OxCJ@xkQ:W6S1bH\\\\{RGGQ3:CED\\\\}G>v.0|5\\\\{34DZ:\\\\{dZhRl@BQgDmBJS0-FxuQINqP--ZQRQvIuvY\\\\{,z6w8zf+ybbBXE/y@VQaybz*30P.7MyJYzTzGUEK,=+eRaqxQ7GBN@U|rTbYH:E1Mz4+G@wOCMFI*b\\\\{b;X,?:yBXleTCd\\\\{PCYaleU@l<ivoz\\\\}b7z6LqRkbOa3LP\\\\{aA23K?YaP*kW\\\\{FUToDi*m10DxY\\\\{C9@<5EcNazbm*7*.bxIxblq?[R39Z0bp:QUP\\\\{py>xg:le//bYS;kbRav"));
$write("%s",("bZVa,JDxPj,ZacG?vtb+|HQj+97<vCUn36bs/GD95yO@x.*KRg>;>n8?aOaybevTOc?ROg\\\\}0bvbxI-*Ta>x716zV<QG0E2x7b5V4W/bL-dT*UZy:Cf*O\\\\}OajxV\\\\{T\\\\{xV=aUat:fBM@;Mwb2*eM2zG;4MIWB>FWAN>?9Iv=+*\\\\}*a*qDU\\\\{j*M2lvQG,?Qa9bzbUa1QRu5.p:-bNawvR64@pyROo\\\\}HUzURvPv/>IS>vTaRaPanRhPybOam-*b-<WKN,S,AzBa\\\\{J-H5DT:=SPJv6AaiFI\\\\}7V5VRa?+WMPV,zm|IU@H3vj/D828i\\\\{*P?4D=\\\\}9/\\\\{Y9?aiI*bmUY-Ga6fFv\\\\{OGaWVSGGByIO6:3RaeIPV-zHV=an3m1s6Sa2bRa9/p=P.j?7vIz7vvbhb0b/Dxv53336/=|p=GS,bUvRuuyL4m.i-:P:\\\\{a;4aeUt,Y\\\\}+NAJNTkbYam.G>@rqEkVGSs;4UGa*zEau6-bVac:py7T>-.b=||bUwNacb-T.b>7<|,?<?.brRNPUaMGu6fzc:4UPaqQi\\\\}6bc:IUwbQdN,S2qy@Ulbd19bdbkvqv>FP*xw6bvb||GGbbP*v/tblb26lb<NjUiFv641LP6b+b1b|54xGam3SajO6bUa*HNaFN7+*H>7t+Bvw->aPw@aJuwb>74akPmTkTt+@al<R1RuEN53HDzw|P*Cax2b8xNafb=a-bJRi5E@K4||XyE@I>O4X<Y*H:JQlEAa"));
$write("%s",("T-2?IQ,b3bzOXCk-Pa=aWa1JhbmEw\\\\}RK;>\\\\}bKRYz>yDScOxbm*\\\\}w\\\\}9eE@QSQ+47HhR6Q\\\\{eONbSPaZRTaj0wbtw-bO;EalbYS>O=Nh4w\\\\}kL?xk|Ca2I71Y,-3A\\\\{R?kQ<SKQ+bL4lxU+m:0vvNbIX-P+yvYaVx\\\\{N|G*wP|\\\\}>H:FDt<ub\\\\}w2bN7WDwPXai.2MB5+Jm+F2iz6OQv*bxvQEu<7b60-\\\\{hSl1TR0Fi..0:9UFLvm+NaV/CCWOMFMMOQ@dMQ\\\\{A2bCah1w2:9w2wzE9mOE,Mtz6ib3y2biFMPWa4\\\\}cHT2.Fh:J<MtPC3wyKd\\\\}|4-,JH\\\\{54\\\\}Evkb<PD8+:@H8b2,*xm+p.EOi1Z83vDzd\\\\}3bzb?x,wmbqz@xSJhFMzIIpI9=wb.4aR+2YQ/*ebiF@aOA@1\\\\}DTPjD2\\\\{KbRGn8m>b462Z?PLXPrgVPS|N<ZeYalb<:m1iQxQHxvQn>pPw;sQbwoxF.V<B.Xxg@wLtvE@OIRGAzXagvDa7vUy:?REYtWym1V<y/M@Wz246Pv;mb>vyvN<5:yODwYaAA3LJ-\\\\{fB,-\\\\{Tzb/HC\\\\{v21R3NKlPxgjPRxl>xLtzb6R+iFRau\\\\}=|B@Ly-Kpy\\\\}NH:m7Q/C@@ajbD/b.wP4\\\\}/0GA<OtK.ChD2PI<Izq7H?ALo-HIaNMHT5NrL4VxXM6Djbj1dM43Bawwm6P/ZO.4,2D?MF=JPNRfNNKxMww:QwOwK"));
$write("%s",("=?E;OO/b|xz5vAwaw2wr+eOQDkC6bb.6>O;6>4>GHMwv8n\\\\},>Hvoxo?K<1w4zb|mwM\\\\}j7hMFFB@*F?@2\\\\}sviMGFr5p@5bE7INfvQvOvMvKvIvpyDa7MU;Fa/c-I4+/yO|6z>7HNkJX-c=>76EJ45v3voCwMuNg\\\\}1v/v-vB+\\\\}v\\\\{vyvwvuvK.4a\\\\}INMEfLMJ=G?\\\\}9DM=|zb<vv|bDl|r0E.\\\\{.tb7+abP*mbi.ibB,9b*b?awwsyvvb-47>E/5v|u5X|pI=LHyw\\\\}JIDJVyxzr+<K/bK\\\\}iJg*DaiFVaOAH/J5H5L?>aEyi/Ey2M\\\\}deFg?BMz?I,BGX>7vz2;H1LG>s5,IjHQL2fOLkblbXah19L\\\\}buwD7M=;MVEFas/twy+GI\\\\{LOa\\\\{b15\\\\{ADaW9K@@DBa>D|6H:|M<xEKo,hLm1?AZ/P*G>PEjIf9i6:KozJ,*bZaT-YFIw@rtbrvuKm=:HW|aBdbz\\\\}Pv\\\\},A?B,3bEa-7SyND4aJFOKcfMKH03wJ8ZwH8>75G-02G5\\\\}*\\\\{-8f<*:ZInx3\\\\{N7U6Qv@H7vhc*@U;RJu*cDwJ\\\\}FN*dIw3kbnLx:zb<\\\\{mG<Co1h\\\\{QB4BXbM:B>B:Sa743:T0zbB/q\\\\{fLMAb6zD2>bKkzxA5>z|NaEav=hbeG1ymb5=q\\\\{AE4a:E>Jre<J?Kb.91M6-,tE|bICK@S0849Jb.tEu5oCOEe9mvMwR10bG@oyJ0T2eb"));
$write("%s",(";6M9*dtyry\\\\{0,GxtXaib2btwz+G4Xyw,tJEA+E\\\\{b*bUaDa\\\\}Elekb|\\\\}M+Wa@8pFR0UaiF66@A20T6mbN/Yu36uyNx2Ef7n\\\\{fFm-xy?a\\\\{3DEl||\\\\}|,E<w\\\\}\\\\}GS3r;b6:1;yvD*Ife|Ihb74m17+ZaKzW/K843N*2bf-abv/mDj+s4/@2|V+EH75Aw<H+FW,GAl427\\\\}9WEx*mvubE@gyNFT1s,O\\\\}7*zbFz4?f:h|X5:FtHW6Mxdbu6|bib58@ac|-cl<.yI\\\\{q\\\\{9>0>a<p,lG1DX5EyN/ivv76b5:gbU7+>R?\\\\}6,.+dR|,bO;GaRyhbn\\\\}.b7+fb4avCkHWgiHQ71A/=Oa79oI\\\\}|@|7+P+X98HJ>R1/\\\\{r+nC/B5?kCyy0y3bv3OHVae<3v|bO4D8Oa4\\\\}1.owZaYaD84;;*@aV\\\\}OeC.|xf<+bP8Oa,xTal04,Oa\\\\}:D0@wXw<7:,xxBDE/6+s|3:I\\\\{jGa|lb3\\\\}WuvEA.GaA**+>**wUas\\\\}-\\\\}B>1A8COaw?oFdHuwZw5:4avBKFOgIFl-@/bbg1?*D.PCN/Y@O;bw/bN*8babWaFa5bvb1=AA<GuGub3bm-P?Ta;,Aa\\\\{xq\\\\{R:I73|iFZa98z@,3*x4AibH3G8eCC.L3J3iFxtLz5\\\\}GaaGn;f21>P4m-x850I;j//ble\\\\}\\\\}0bleny7vxbCDp<*4Va=|1C>5B,XC85w:Oan3|bT7EaG=Z@O"));
$write("%s",("vXaCCbFt4E.U<RvH|4akA;E-h9ET1D@*FP17/C7?aNaCv-bZa7b062xdE/A3\\\\{tw5bhbW/xv5w::kb7bwv*bu5s5fbK2RDjb|\\\\}UaW*0bbb,,0b7\\\\}5\\\\}c\\\\}u8.bTyJD/:H8/bfDdb+9d2fC|9*,R@x.M7G;W6=-a7k-<*.bF37b8?6?EvQz+dTaI4\\\\}9N\\\\{\\\\{bf:3:tbE@:>/Cy;g5i74aW?wDThuD@amEvbr@I3*@9DeDkb@AR/xAR-xwibN/sw4vcvXbcvKD\\\\}B2=Ra2b.CNa?aibubYaibzbkbVaS@w1uwt:FB>a:4Z2swA.Pv\\\\{yP.8vuAz;le.b5\\\\}czX/cb-+1,/babI\\\\{m1uw8.Ea*|*AZ31vB,|7I\\\\{ib@xr>Iz,zI/l1Xa.+f-J+\\\\{b3yibi/UAMAdbk\\\\{/xRBC?Xa4aS>wCyhuC5bg?w?Gar?5;mb3\\\\}KCh\\\\{\\\\}25Bk@lBQADa\\\\{@d@jbR,@a@wf8C4EBVy*bs|=a*+wbI*L?Vv>56xOxg,Z2<\\\\}w2w=2/*b2/QaT6-bG;79\\\\}AYzYa0=EB:4t\\\\{y?kwUA,@p?:8N>/b?8lbmB0+=>7>bbb.4aX=wBDguBE@L>Oamb\\\\}wd?7?b?DaQz?aNB@a>7F82bm:UaD.Sa8b309BMt0x3bK=FA,4s7348>m:g>YaSaRambX5gBd;,bO6t\\\\{Pdz3,5C-85X9Xb,:b95b2bF0zBIxI?E?owvb>aGa:cXw2=p=97gAC="));
$write("%s",("H*\\\\}94a7<lAshjAn3XA>ab.Pa46d\\\\}H:+@Paxbdbo8m80APw:3c6a<f?Gak<z5jdMwg/L49b7z\\\\}@\\\\};6--@S854Qas5p136a-n=h>/:XajbO>88F79-tbwb-bcv5:\\\\{+o\\\\}1wwyDa4.I|O@k8Pa/bmw?<y+Z;q1Pu15@5czy@-+G9,bi/s@VvO,5bM8:<=9X?phV?2,S46;<@:@9.\\\\}\\\\}\\\\{4Oahxzb!![2iba!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"o3j[2|pa\\\\})3(f\\\\{#(tnirP;)R3FZ0=af+=awb20XbA,Aao8e;A<0bhbo<M7\\\\}9pw9,ovi>g-;\\\\}hb.b7\\\\}H3lbmbdv0b\\\\{b-bcbbv?*K-abj,3\\\\}d1O*hxH:S/cz+wW;q>K<24j@\"\"),\"& VbLf &\"(\"\"L4Z5>aw1hb*dM,>-<-V-Dxg9g@r7e@q?Bxubk>93T3p7Q<b/U.4ab8T>VgR>vzT23bTaPv7b23|+5blb,bHz/-04abebm>m2,=y06btbzxlbY\\\\{yb<vFa0vi9dbg92bVaQz3b03,b6,gzlbjbM:R\\\\}E+b6</s\\\\}V7M=Z2i|Rz+e9=H:Dxz0+bf-y*Va.2lbL4x,,/L=pxIzh9"));
$write("%s",("+eZaQzH:uvk6;\\\\{H6Y=-gW=y7Pze.8>G>fb\\\\}9m:m1i5P.+bVaz0Z<XaU\\\\}4v2vK-N<ixd=2>98P;k08b3bB+jbS:?+*9w8Jz-\\\\}4vI4wyYa3bVa9/AaPyRaOac>@aNxV;T;1yA2l\\\\{-4w\\\\{a4W1J=Px2bez@tWaTaZz4ac58<Li6<>4y:O=Wa2==4R1Vay=W9,=w,x;92Waz:K-SaEa/bh;=aEa4wQas6Vam1\\\\}9n3*=h;p=WaEaSaVagbB<q:N-hb.;0\\\\}j4u=Aa.bRaEaabVaTaVa3bo+@amblbM\\\\}J9x7uw\\\\};/bTaY\\\\}t4fvI|D9-blzuyOaN+lbib>aww/09z1-abh:f:m1P:81kb4,Wazy,bf-Va3:o8s:c;f\\\\{Y;K-bb@,:94aO3>92i<9ebG9ybAaifG*bbQjN+.bk1u+Q.38z;cb?:M;9xabhxv:twNay+/;69F-,\\\\{le8b<;gb3:K*8beb0b>vX90;F;@:Nxub<a,bjvhb?a24Q:jbSa4+Da\\\\}bSaK5z+,/V9R9p\\\\{tb.*x.h10vh+7bAay/mwh+0vH1F1wb.bdb<a<\\\\{r++/n:j0g:/:B9kbD.9\\\\}mba-y7l:vbk;2\\\\}eb5bNav73:Xac\\\\{|7gzMtTaUawyt:Awr:Fz:yUt:yQt:3:9W8G.zwB1+9c.|8v.dvvbc2Oa5:;8J7U7@aNa+6Vu<a\\\\}9T9?\\\\{dbQjQvbvQvrw1,Ea3bBaYu=aSyV-axtb7bW08bm"));
$write("%s",("bYaU\\\\}xvVa8bWaG9/bAa3xn8l8*bjbNaf\\\\{U9P.vbf8Z/8bAaTaFa+bFvZalxRawbDa>a89o,|9bw\\\\}959kbL\\\\{29-b=alb@637+-,7Da,,o8G|axm-E.u-p2c8ija8ab8b<\\\\{X6xz|2Ra:.h+vxz2Ww-b+bQv:86-B6U4ubr|K3qw,.mv4\\\\}tbmb;6+b@a>a\\\\}.lbPaAz9.r+Qum8le0bg\\\\}Eawbd\\\\}kbib<xy-00wygvf/ybNa@av|x*Kz80y-hx\\\\}b*1Na=|kbs\\\\{cbk+i+g+Va-+r\\\\}D,3yjbJ/u*67z|y1t1Qd|-Ty6/RaK*C7CaXa.7y/<vZap\\\\}Xa6vNvLv7bhx6bVaIw/b|.2xdb>aJ5Z\\\\{:4xzn,Pu754aM0I6xjG615@a,bDam1=a15/0z1d/wz.0cbkbp0K/C6|1Vy/0e/n\\\\}-b\\\\{bubu6ebo+>au5=\\\\}lbcb7bR4tx5-K.j6T1h68rXa\\\\{bD.++Xar|C,y*mbtbM\\\\}?6+xf-Xaq5=1:3Hz83Kz9-m14-l6@6Y0k4J28|g|,6*64b\\\\{bL42b2*V|:3\\\\{w/b7/kb+b>aNa0b@ad\\\\}yb4aX.d5Uib5vb1bf.W4=\\\\{Q.V1i6F|@aXaQa4bDaC03yUaz6\\\\{bjbfbCvUaZa7||3+b2bd\\\\{0bDaf|8b7+6/HvUaEaEaAa80\\\\{b/bWag/R/\\\\{0w,Z-X-I.wyt5Sac|Q.U4h/Aa,3gb2/Ra?\\\\{cbHz.5Wa,581"));
$write("%s",("Iw=am+DaubWaif-+tw8b|vdbC-75Ta2vWaC.mbl/j/>a25Ew?v\\\\}\\\\}@aDa?w@w6bAaY3JwWa|b<aV\\\\}lbAa5,D+tw1bib=,cb<\\\\}nzx*8+CaY3avD\\\\},x9xmbM\\\\}U1a/r-P3OiN3hytxI\\\\{w\\\\}e2rxw49.0vG1lx73Uafb\\\\{0P.\\\\}\\\\{7v\\\\{bj+8.+b9-?-b|/0RaVa\\\\{dSa?alzNa,bhbCaZaK1-bEaB2tx@2c3d4Tz?1b3f\\\\{k2vbD0y/5\\\\}\\\\}w<\\\\{r13v2\\\\}s|*bN/Vwwb?aH2Z+u,S1Va/bfba|=3\\\\}bdbc3h\\\\{V3Mv2b*+*2<142A2224a;+q2Kio2h+ibBayy/b4\\\\}yvf+yvN+4b*b6x2b+bkbQah\\\\{a352Hx328+wv\\\\}bab0b|*AawvVa7b>aUaUaibUaOa2b=a0b@|lb0y+b6b,bB.Syryuble1bqw|-6bjbn.SaMvvbCz>2*2u\\\\{*/tz,vY\\\\}Na9.zb/bBafbq/1bUaybQ1vb?acbz2y\\\\}8b6b-bHz51lx31Tzx\\\\{?w8|Oa.,yxkz*2=xe\\\\{Wz41b+DatbxvVyy\\\\{t2>17zl2;1Bcib:wgcYaVw21T14aG\\\\}N0FiL0,x=1o,w+5vF,Qj*wq\\\\{A1>|3vxy6xi0fbj,rvv,Y-Rx01lb;\\\\}.bx1v11bt12bkbcbGzPaEx7bUaA+d+I/.-11i\\\\{v\\\\{t\\\\{CaNa|b@a-bHxFzt*Dzk\\\\{X-X+evcvizu"));
$write("%s",("yabB+m1JvUa5b:-cb\\\\{bibuz6b2*x+ozlbx*jbT/Aaz0E.NukbAanzz+N+Bawbg.QySxAyRa7b?ePa.bS,xb4a8\\\\{Y.uiW.Ea0bUa8bCxRa-+Bale\\\\{fP\\\\{7|B+\\\\{b|\\\\}Sa4bhbWaUaz+\\\\{.Uawbkbo+m+PvWaCah+/b@awwmwcza0gbibdbQvjbD.*xmbK*kw,bPaTaAambgbmb|.Hv7bcw?-=-4-2-jbXaKzWa.+uwK/\\\\{/lzabcbAa/bXaXax*zw@+d.G,c\\\\}zbB+zb+bm-V,1bTambj+Zzeb?aS-7+Pa4b@a4\\\\}3,\\\\{vh.c\\\\}=|8bWvq,U|T.XaVxH,\\\\},ibJwuyEaB+O-1bY,/b9.5bL\\\\{-+dv,b=aCawwzbz|DxTa6zNx4a8ys-ciq-2bxzS|F.XyDaJ.C-d\\\\}s.jbrvh-bb\\\\{bg.kb3bCaab1v0bi\\\\}hb6wfvOykbb.cbtbib6wib/bSyFaN->v<a/\\\\{.\\\\}MzM,K*D,XaebjbAaBaI-Rar\\\\}\\\\{f.bn.o\\\\{C-?v*b2bf+bzd\\\\}*bO|FaVx7-t*jxuba-L\\\\}?a,--,Wa?afbhb3b4\\\\}FaOa/bcbQj>aeb|bmb*dbb7+.+=ai,WuE+L,XaAa\\\\{bc->aTaw\\\\}v*lxs*AaabDx,bHxVzy\\\\{@zt,Y,wbIv\\\\}b4yq\\\\}Saf+wbj+4aiw<+pk:+Za-bixZa,bSambw,Z,=\\\\}0bZzlzjzsvS+Y+8bixmz2bN+UyQv"));
$write("%s",("=\\\\}>aLwx*vbVa,bZzx*w\\\\}1+m+fbib+bBadb-b|\\\\}E+XwEatx0bb|zbf+ywlbgb-bSatbcbvwCafbmb3bB\\\\}n+MvQ\\\\}\\\\{xjbbxDa5wR+K\\\\}-x>zxx1*yzT|e,bv7v.bizc\\\\}+wMxt\\\\{Zu\\\\{fifDyubM\\\\}Q+7bQyEay*k\\\\}+wi\\\\}g\\\\}zbqwcbjb3bi+ibhbtwOe3vvbSaubgbVxv\\\\}n\\\\{4afwH\\\\}kkF\\\\}kx/bkbSalbO*Faq\\\\{c+abdv8bOaMvXuK*5z3y8bEa|zq+R|Ca=|5b2*5\\\\{0*B\\\\}Sa3bYa*xEa1bab\\\\}bNvdbw\\\\}p\\\\{u\\\\}8rSaP*N*|b6bkbFa?aJvRalb*b/bPa1xBaebXv+y8bJwl|izl|Oa+z\\\\{bJwLvmb1bVavbdbBxmv.b/yC\\\\}fbE|*|\\\\{z3\\\\{*w,b6bWw4bmb6x|bZaK|\\\\{b.\\\\}q\\\\{o\\\\{vbm\\\\{t\\\\}V\\\\}uvV\\\\{yblbTa3\\\\}vbjbRaDxVv\\\\}bhb,bTa|bNapw4b+bTaZazb6|fzkbWa8zubDaj\\\\}h\\\\}/x4aWt9\\\\{3k7\\\\{Qx,wubVaybVbdbcbWa.bb|FyDypwZa/btbgb.bAaTzPas\\\\}Da8bhbSy\\\\}bmbBaVw,vQajbkyNzLz\\\\{b1bdb8b.bTaQaOaXyrvNx-b@aQzbzkbgb|b|vzvxvvvDa|z4\\\\{mwwzs\\\\{QaTa\\\\{bUa\\\\}wab>av|ixgbnwQzybDa.bow0\\\\{,e@\\\\"));
$write("%s",("{>\\\\{Saqx9b.b?aebzbNahz;zVa5bRatbr!![2iba!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"o3j[2|pa\\\\})3(f\\\\{#(tnirP;)R3FZ0|+wYatbRa>awxlvv|lzSamvAaEadbSaBacbmbmbXa>zoxcb\\\\}b.b*w/bVakbNaxbevfbkb*bTaNa5b?\\\\{levb,zGa.\\\\{tvcb:vLw3bVuvw0bPa,wMvybRapwAzMwle3b,bvvEaqx4aSt9yGk7y0v,bzzt\\\\{uz\\\\}\\\\{Cale-b3bUaGa9wRa0b/yebBzj\\\\{vdg\\\\{hbKxYa\\\\{wOzNaMztxRuUzSzQzub@x>xxzvzFaebOaozmb\\\\{bIzGzEzCzgbAz?a?zzwUx;dNaExib,bEa7bGxOaExebTa2xRaSxhy5bizgzezSa5b.b?x|b7b-bFa>a+bjbUavbzblbleebWvpxEv+bhb<xlbJxQazbUwRazb;wXaSa\\\\{bWaVaDxubQa\\\\{b.bUaab5b<aOy|b\\\\{bkbdbvbOatble*b@aUaQaPawyuyhb>a*xmy<wMv/b=a1bPw4y2y-bDvdb0b4aRrgw;khwPwib0bZayxUaPa7bDa*d1bWaVvzbAatbebmbibTadbmb.b-bdblbyw"));
$write("%s",("*xab3vzw3x1x/xQxfvhxZxBacxaxhb*bXaEajb4x2x0xFa.x,x|b/b?x2bmw;x1bEa0v>amxsxOaYaEavdYaFa.bmwabGv+v3bAa0bdbzwWagbwbVa?aLwSa,bfbcbiblwbxbb|bDaqx7boxmxZakxWvYa0vTaOavbSuAv3bXabbhbNaBaDa1vtbabubhbTaab.bmbwvBbjbPa,bAaCaFatbWaBaabwb*b+vPujble?wDahb7wgbvbNa1ble7b<a>adb/bSaXaFagb,w-w+w\\\\}w/bYagb7bxwjb*bAaFambSaYabb,beb1bfbwbhbjbcvAaSrukewTtXjVtXacbhbRaubcvEa>aFamvkvfvXaabzbEaCaeb-b/b-beblbzb,bNa7bvbkv5bJbPawb2bBajvlvgvQdZamb=aYaab,b7bmbdb.bOaCaDa|bEaYaeb.bWatbdb5bmbjbDadb+bmbDa7bNaCaEazb2bRuvb2b0bcbwbSa1bZa|bWaubab7bZaBaEahb<aCabb*b7b?aQaUs4u2s.tEt5ueurtiubuUrJsmu3uyeou+u;aVr:tItPsNsXscu|tsujuyunuwu-bUsttCatsFtguDtwbWbUs+tusxg/thuPafuEa@aXsLsjt@d=tBstsktUs;s9s/bSrokRt9aSr=jQr-b4bye\\\\}fubjdVrot,t2tlt;t>t9trs9aEaOaJsrg3t*tpt4thtZd:a-bJsxgnt=aYsRfqt?sctuths2sVs+sTs@a<"));
$write("%s",("a-bVrRs4satYsEfWs0sitbt|sWezsJsRfHsZs:aCaasIsQs>aAa-a2fssKsxs\\\\}sms=sDsAa?a>ats@sbs>sEf<szbis5s*sFaBaWe1sysls2f.s*bvbtbRe?fVr/sjsvsyedsqsFrosOaVrpsws?aAayersVrZris\\\\{d-acfescsasksYr9aasHareOr8aCa@aWe*f\\\\{bvb8aUr0e8arb8a8a2b4a4a+j4a4exb3bCb6byeDbbcubHacfDhfeFh3b4b.b4eQbye,bMbKbBb?ahehoYqurxr.r0r\\\\}rgr\\\\{r|ryrzrqrwrYqorvrsrTqfrprmrrrkrnrhrSqdrerlrirjrarcrZqCqXqOqbrMqVqWqPq@qRqIqUqQqGq>qNqvqKq6qLq3qHqJqFq\\\\{qoqEq4qDqAqBq?q7q<q=q:q5q;q8q9q.q0q-q1q2qwq,qzq/qxq*q+q|qyqiq\\\\}qXpqqtquqrqsqhqpqmqjqkqYpbqlqnqgqKpeqfqcqdqUpaqCpSpZpWp>pJpTpQpVpOpRpLp=pHpIpPpMpNpEpGpDp-pBp9pFp7p@pAp:p*p<p3p?p;p1p|p8pZo5ptp6pqp2p4p0pepSo/prp.p+p,p\\\\}pupzp\\\\{pxpspypvpwplpnpkpopppapjpdpmpbphpipfpcpMogpBoUoXoYoVoWoLoToQoNoOoCoFoPoRoKo5oIoJoGoHo?oEo-o=oDoAo|o4o>o;o@o9o<o6o\\\\{o2o3o:o7o8o/o1o"));
$write("%s",(".ofo,owo0ouo*o+oxoaozoqo\\\\}oyoooYnvomosoVntoNnporonoDn:ncodo=nEetbOjEg>lGmeoZnOnboWnTnXnRnUnJnLnMnSnPnQnFnKn/nInCnGnHnEnBn6n@nAn>n7n<n,n2n?n\\\\{n+n;n8n5n9n.nqn3n4n1n-nxn0nvn\\\\}nzn*ndn|nanpnyntnwnrnZmnnunlnonsnmnenJmcnVmjnknhnTminfngnXmbnWmEmYmMmOmCmUmPmRm@mSm8mLmQmNm\\\\{mKmHm.mxmGmImDm9mFmAm>mBm<m?m4m6m7m=m:m;m0m5mmm3m-m1m2m/m,mtm*m+m|mumzmjmpm\\\\}memimymvmsmwmlmUlqmrmomkmbmnmZlgmdmhmHlfmElTlcmXlamVl;lRlYlPlSlWlQlIl+lGl7lNlOlLl5lMlJlKl9lFl8lDl:l1l<l\\\\}lBhre3e<iHgMjbl/lzl6lbl3ltl4lql0l2l.lglTk-lrl,lul*l\\\\{l|lylvlxlnlwlilslmlolplclllfljlklhlZkdlXkYkVkelalOkPkMkUkRkJkNkWkIkCkQkSkLk3kFkKk@kEkHkBkGkDk?k<k+k:kAk>k,k2k;k8k9k=k7k4kyk0k1k6k/k5k-kvkik*kuk.ksk|k\\\\}kzkgkxkok\\\\{kwkmkdktk=jqkakrkXjnkpklkBj3jkkYjjkbkhkekfkKjckEjZjJjGjHj>jIjBi|b|bvb?e.b3b>b9dLg:iRfFjCj@jAj9"));
$write("%s",("j?jDj8j5j;j<j.j:j,j4j1j\\\\}j/j7j-j6jzjqj0j2j+jijwj*j\\\\{j|jyjpjxjujvjsjtjjjajnjojljmjrjkjbjhjUifjgjdjejVi8iZiOiXiYicjWiHi6iTiKiRiSiPi0iNiFiQiIiMi-iJiLiGi|iEiuiDi3iCiki2iziIhzbDb\\\\}frbZdlgKgYg2i7i4i5i*i/ivi1i.i+i,i\\\\}ixi\\\\{ioiwimisiyiqitifiridiliiiaipiYhginieiMhhijici-hShbiWhZhUhLhThQhXhOhRhVhPh.h\\\\}hJhKh8hNh6h9h*h,hyh:hpg2b3bSeHepfRfmf2fkfJcWeyf-bDg3hwh7h4h5h2h/h1h\\\\{h0huh+hzhMg|hshohKgxhphthGgvhDgrhVgqh:gmhWgnhUg8gSgKa\\\\{b;a.cwbldIaXbVbTb0a9dBgigPaPgTgQg6gRg-gOgEgNgHgLgIgJgAgFg@gBgCg.g?g9g=g>g;g+g3g<gzg*g4g7g2g5g0g,gwg1gYf/gfg|gyg\\\\}grg\\\\{gcgqgxgugvgsgbgdgggtgjgSfTdag4eybEbCbXd7dXf1fcfegWfZfUf;etcQfRfOfVfMfPfTfNfFf?dDfEfKfLfIfCfJfGfHf-f/f3fnfBf2f.flfGe2e1atc1aobwcubwble,b9dIdge6e9efecf,fre+ffe1bldwb+byeZdVb8b1bEbxb;a:bfe6a@d1d5ecfqemcZaWeQehc5bAd:eVe-ctbld"));
$write("%s",("-are0dFcDc/byewbwe3bxb,b;a<bfe:breaeye8bEc,bxb2b2btb;a?aWd7e>dmereoe7dpdfeEbYdHafe-e-eFaGakexb-bFc4a-afe.b\\\\{b+cMajaPanePcfe@dIdeeGa+bxd9dSdPabeGa5a@dSd3bDbBb9d>dHd@dobIdRaYaOaVafbVaib9dob>d6d4d-a?a;a>a-aPaBaxc7dVaNaUa?a?a1d1d-aebcb/a1dxcvbpbEaVc7b@aFa@aAa@anb+btbub.b+bzb>bMaHbNc5a1b3b2bDc2b>b:bpbDaBaBa;a;a=anb-bVc|b-a!![2iba!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"o3j[2|pa\\\\})3(f\\\\{#(tnirP;)R3F#cWbybHa/axc-bxcGb:aIaDblc:avb|b+bub4bcb-b.c,c*cHaQbJaGaxbNb-b8a1bxbwbtbxbUa-b.b|b3bvbxbfbucsc3bHaHbtcsb/atcobJaub:b6a5aDbtb,b-awb|b.bibHa7bxbzbxbeb-a3b1b.b/b,b|bHaebdb-a,btb1bzb.b1bAbob5a3b-b|b1b/b/a5aJa2bm6Aka721(f\\\\{#,43b7Bja8361(f\\\\{# D4[O31da172Q"));
$write("%s",("3a3:[R34ma5114(f\\\\{#q\\\\})4;6c:6[F52da49996[E4:ca46j:[O;?ba&[2iha=s,y=z,Y4[O32da827-8[R38ea9909-8[-8?haq\\\\})2594:6[C?9da3418?[YD[D4[YDtca42t8[XD:ca939?o=6[\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'8[O3~07[-6:ba01?Uea0804wL[G5;27Gi:[D4[;F-ba5[BGt8Oda874lLoyay,]99999[gnirtS wen=][c n3aea\\\\{)v]y3b&a(niam diov citats cilbup\\\\{RQ ssalc17[w9[D4[w9oca38v9[v9:ca97GW[(ICca0696[(I:ba3TDaj:[HWB8a cdln&&&&;maertStnirP/oi/avajL tuo/metsyS/gnal/avaj2>b&ategn&&&&2 kcats timil.n&&&&]; V);o?a;3ecaL[\\\\{?av?hha dohtem;3a/4nga repus~3acaRQ83cgassalc.X6[-:2ca30%L[-::ca53!$Ka-:[M?4ba0B?G06Nda9928A[M4Bca57wVa96[;56ca62j:[8ABoa(=:s;0=:c=:i;),@ajaerudecorph5[hY3ba0iQ[R3;da63588[ZYBda886-N[N?;ca67C?[AS[D4[O3rca02gP[s8:ca71gPara&(tnirp.biL.ok\"\"),\"& VbLf &\"(\"\"en\\\\{D?bianoitcnuf6Y[O8[D4[XJ*ca23O8[h>:ba0iIaYJ["));
$write("%s",("YJ?ba996[95:ca45j:[|[9ba0D4a06[!$W5tPbqa(rtStup=niam\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'tni5L[5?=kawohsn\\\\})291jIFi<Mca1488[:5:ba2<5a.6[YQ3ca28i<[;5:da454/6[;57ca099?[?=<ga4(f\\\\{#=DF[-A>~?b%a(amirpmi oicDAx\\\\})6904(f\\\\{#3Cx\\\\})633Y[3Y<va92(f\\\\{#ni;RQ omtiroglag7[\\\\}G2I6bL5aea.tmf/Rcfacnuf;Y4[Y49datmfE4[E4:raropmi;niam egakca|I[lB4ca02?8dbap/8[I4:ba-C4[C49jatnirp tesK4[xI3ba0:Paban/P[VC7*a15(f\\\\{#(,s(llAetirW;)(resUtxeTtuptuO=:P6[p>3ba5@8fG4[G48daS CE4[O39ca&(C4[.68ba x8[x8[E4[O3\\\\{iaRQ margo76[O3;jaS D : ; R>6[O3:ba\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'C4[O39qa. EPYT B C : ; AR4[;6:ka)*,*(ETIRWM4[E6;haA B : ;K4[O39ba [2cJ4[;6<ba:G4Is[Cga(f\\\\{#(>\\\\{MBba3hOabafiOFba5aPa\\\\{aetirwf:oin\\\\})8(f\\\\{#>-)_(niamp3cL6Bka(f\\\\{# cnirpPIBb6a,atnirP\\\\{)(niaM diov\\\\{noitacilppA:RQ ssalc[\\\\{7B%6ew4aram diov;oidt"));
$write("%s",("s.dts d[ar4?kaenil-etirw~6|va(,\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'s%\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'(gol.elosnoc;)\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'x4/[2kya\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\' nioj.)1+n(yarrA>-)n(=f:4\\\\{ia!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\}54,1\\\\{.v3kka# qes-er()y3kba&)6.ba!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"E3lD3/#3.h40la1% ecalper.-6|@3k6Bosarts(# pam(]YALPSID/8kua!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\".NOISIVID ERUDECORP&4\\\\{ma.RQ .DI-MARG23#j4do"));
$write("%s",("aNOITACIFITNEDI+3kra[tac-yzal(s[qesodX5c\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'a!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\")!!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\");\\\\}\\\\}!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\");\\\\}!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\");return 0;\\\\}/****/e3a\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\");s=\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\';while 0<len(d):\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\n x as int,y as int=d;i=3;if(n=(x-5)%92+(y-5)%92*87)>3999:\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\n  for _ in range(((d[2]cast int-5)%92+6)):s+=s[len(s)+4000-n]\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\n else:s+=d[2:i=n+2]\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\n d=d[i:]\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\na=0;for i in range(len(s)):b as int=s[i];a-=b;print((\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'+\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'*-a if 0>a else\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("'-\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'*a)+\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'.\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\');a=b\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\");gsub(/!/,\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\",s);for(print\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"define void f(n)\\\\{\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"00g,\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";for(m=128;m;m/=2)\\\\{\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"00g,4,:\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";if(n/m%2<1)\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"4+\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\",\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";\\\\};\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"4,:,\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\}\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"389**6+44*6+00p29*,\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";++j<=length(s);print\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"f(\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"n\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\");\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\")for(n=9;substr(s,j,"));
$write("%s",("1)!=sprintf(\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"%c\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\",++n););print\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"4,:,@\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\nquit\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\}\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\")');\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";FORiTO UPBtDO INTn:=ABSt[i];print(REPR(50+n%64)+c+REPR(50+n%8MOD8)+c+REPR(50+nMOD8)+b+\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"J\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"+a)OD\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\"\");end;\\\"\")\\nsys.exit 0}\"\")]]></xsl:template></xsl:stylesheet>\":s=\"   \":For i=0To 7:s &=Chr(32-(Asc(c)>>7-i And 1)*23):Next:System.Console.Write(s &n &Chr(9)&n &\"  \"):Next:System.Console.Write(n &n &n):End Sub:End Module"));
end endmodule