module QR;initial begin $write("%s",("Module QR:Sub Main():Dim s,n,i,c As Object:n=Chr(10):For Each c in\"<?xml version='1.0'?><?xml-stylesheet type='text/xsl'href='QR.xslt'?><xsl:stylesheet version='1.0' xmlns:xsl='http://www.w3.org/1999/XSL/Transform'><xsl:output method='text'/><xsl:template match='/'><![CDATA[write,format=\"\"%s%s%s%s\"\",\"& VbLf &\"(\"\"\\\\write{-}{txt}{(\\\"\"with Ada.Text_Io;procedure qr is begin Ada.Text_Io.Put_Line(\\\\\\\\\\\"\"print\\\\\\\\\\\"\"\\\\\\\\\\\"\"STRINGz:=REPR226+REPR153,a:=z+REPR166,b:=a+\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"2\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"+z+REPR160,c:=b+\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"8\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"+z+REPR165,t:=\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"write('implement main0()=print(\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"BEGIN\\\\{s=(\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"#include<stdio.h>\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\nchar*p=(\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"Ra#include<iostream>!nint main()\\\\{std::cout<<(!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"class Program\\\\{public static void M83apbSystem.Console.Write(!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"let f(c :Int):Latin1=if c=127then!!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"!!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"else(string_of c@!!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\" g caffeine !!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"@$3kEa!!!!n!!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\")@f(c+1)in print(!!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"Quine Relay Coffee.!!!!n!!!!nIngredientsq3aha!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"@f 10U3cgaMethodz3c#a);let g(String ->[])!!!!n[c;t]->w4edaPutY4spa(int_of_char c)05auainto the mixing bowl|4ejag t!!!!n|_ k4gtaLiquify contents ofE3oeaPour\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'3w\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'4elabaking dishv6biaServes 164doain g(!!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\")))s!![2aca!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\" [2bo3cparts(nltnirp(])]v3cja.NUR POTSp3cx3dp3jba!!M3dp3df4fda[))j3ci3e,3cp3l[2kga\\\\};)06xu3n<3|pa)1(f\\\\{#qp]\\\\}\\\\};)0,33&*3&+4\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'*3\\\\}ba3R3RA5Mfa(f;)1>6Nba.G5[G5Dba3+9[F5[F57ba7F5NE5[E5[E5[E5[E5[*3o1DlF5[F53ba418[N4D$FOGA[.9FkaD ; EYB RC99[%<[W38da,43H5[H5[W37daDNE78[I5[78[H5[H5[MOtca As>[L5[:8[H5[H5[*3veaPOTS88[J5[88[H5[H5[t>ws>[K5[98[H5[H5[*3toaRQ margorp dneB8[T5[B8[H5[H5[*3sbaS\\\\{>[I5[78[H5[H5[*3[E5[38[H5[H5<ca5148[F5[48[48[H5[48[*3fba&@C[68[68[H5[68[zIvgaPOOL R$I[>8[>8[H5[H5[*3tea\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'&"));
$write("%s",(",)88[J5[88[H5[H5[*3sia. . TNUOw>[O5[=8[H5[H5[W3uearahc6I[L5[:8[H5[H5[y>vhaB OD 0 z>[P5[>8[H5[H5[LTuS3IG5[58[H5[LT[X3*ca)ANC[88[88[H5[88[*Zw%Z[98[98[H5[H5[*3uqaEUNITNOC      01D8[V5[D8[H5[H5[sOu\\\\}>[I5[78[H5[H5[lOv5I[J5[88[H5[H5[4Izba.:8[L5[:8[H5[H5[H5tja1=I 01 OD>8[P5[>8[H5[H5[0IueaA PU;8[M5[;8[H5[H5[*3[E5[38[H5[H5;ca51I5Nxa;TIUQ;)s(maertSesolC;))b6[K8[K8[H5[H5~ca13I5NbanP4Qba2P4O+:[+:[+:[H5[H5#ca3658[G5[58[58[H5[H5sba2OEOca\\\\};88[88[88[H5[,K$ca52J5Ndamif:8[:8[:8[H5[wK%ca15>V[G5[58[58[H5[q>[*3gba+n>[78[78[H5[78[*3u%a315133A71/129@31916G21661421553/l6[U8[U8[H5[U8[Y3ueat+s+L5[:8[:8[H5[:8[*3[G5[58[H5[\\\\{O[Y32oaamirpmi oicDAxd5Qba6qFQbaCS4Rda1213<[P4Dba0N4[y@Eba3D6Opani;RQ omtirogla>=[,@[,@[H5[cF[>Kv~anirP.F;\\\\})1+69%%))n(tni-i+512(v4IU8[U8[H5[U8[Y3+bawH5[68["));
$write("%s",("68[H5[68[1>vhaaepeR.SvW[?8[?8[H5[?8[*3ubaWH5[68[68[H5[68[*3tfa=+s\\\\{)L5[:8[:8[H5[:8[*3t68[68[68[H5[H5#da11568[H5[68[68[H5[H5rea3201K5Nda\\\\}\\\\};:8[:8[:8[H5[H5#da844J5NP4Qba0N4[N4Dda995$<Odadne%<[%<[%<[H5[;8%ca02qMO&<[\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'4[N4;da688&<OnaPUEVIGESAELPnc5Rca29c5OI8[\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'4[N4<ca714<Oja1,TUODAERL8a1?[\\\\{B[\\\\{B[H5[AK#ca260<[0<[\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'4[390ca640<O~a(etirw;\\\\};u=:c;))652%%)u-c((||P9[><[><[H5[H5#ca13><[><[\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'4[)@0ca77><Oda#-<69[$<[$<[H5[H5~da230$<[$<[\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'4[N4/ea3603Q4Nda||iGE[&<[&<[H5[H5$ca54J5O%<[\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'4[N4<ca53%<Oia#BUS1,OD:9[(<[(<[H5[(<#ca544:[(<[\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'4[N4/ca46(<OOXbia)3/4%%i(e5Rba7:K[J8[\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'4[4<0ca28J8OE6[\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'4[N4;ba1kSPba)iC[RE[RE[H5[68#ca17\\\\}<[\\\\}<[\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'4[N4/ba4g@PgaESAELP89[&<[&<[H5[H5~da324&<[&<[\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'4[N4/da276zOUQa\\\\}2=:/t;2%%t+2*u=:u\\\\{od7 ot0 yreve;i-=:u;1=:+i\\\\{od))1(evom(dro=:t elihw?s;)s*||.:[x=[x=[H5[H5~da850x=[x=[\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'4[390ba3cPPha#-<1,OD:9[(<[(<[H5[H5~ea96724:[(<[\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'4[N4.da623(<OBFb3Y[)<[)<[H5[)<$ca74)<[)<[\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'4[)<0ca16)<Oban1KRca02=8[=8[\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'4[E60ca88=8Oladohtem dne.H8Rda529b5OH8[\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'4[N4;da1713<OganruterC8Rca74)@PC8[\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'4[VG<ba4VGPCaV);gnirtS/gnal/avajL(nltnirp/maertStnirP/oi/avaj lautrivekovni$9Rca31uPP$9[\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'4[E6<ba8FW[jQ[SS[SS[H5[*:tca30\\\\}<[\\\\}<[\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'4[rL1ca83Q4[E6[\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'4[>W/ca33E6Oeb\\\\}\\\\}\\\\}\\\\};0=q;)]q[c=z(tnirp.tuo.metsyS;)0(tArahc.y+z=]++n[c;y:"));
$write("%s",("]q[c?n<q=y\\\\{)0>2%%++i(fi;48%%)31-)i:3c&as(+87*q=q\\\\{);07951<i;(rof;n)rahc(+K>[9A[9A[H5[N=#ba4M=[M=[\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'4[8A[*3[E6[*3[E6[E6[\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'4[E6[Q4[E6[*3[E6[E6[\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'4[N4Cca837HO4H[~K[~K[H5[|<#ca70|<[|<[\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'4[g@[*3[E6[*3[E6[E6[\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'4[E6[Q4[E6[*3[N4lea3381Q4N)a=]n[c);621<n++;(rof;0=q,0=n,0=i tni;tE[bH[bH[H5[H5~da449Z8OE<[\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'4[0@[Q4[E6[*3[E6[Q4[E6[E6[*4[E6[*3[bByda692Q4N,b6aeeicpbocLhLf7m6ghF6g2?\\\\}bJaMa\\\\}bJaPawb-e-bJaJao<JaJaTaJa8b<n;a8bSaTaKa8bSar<Tawb|0PaOaSaSa7m9bKa8bWQ?ar<>+Sar<7m+BJaLaJa8b>+7mr4c\\\\}a8bNau67m:b2?:Y2?:Y|0JaHaJa8b73akaHaJaJaQai,~4a=bUa:aUa:a<nocXbddxepgXcVcScQc/aDg|bCtIcncDcbj@c|bKa<c=a0c@aEa2a;c9c7c6c4cAaGa?ay:Ja|bxekcpbzc-bCdlepbocHazcHapb6a6aIc7e=a-ayjed3bHd6a6a=a-a?aF.9"));
$write("%s",("i3fdb:e7apbVRFeDeBe@e9apbGeEeCeAejd1b;.Yb|dCbqi<k7aVR/h-hMayjedvfvbJa>a2a,g*g*hMa?aF.CfXbybvd6a13i4bHdtbq;vdie=aSeRa\\\\}Obf\\\\}O5mgbXaNaSeXhqe7bRhjcYcWc6aSdwdeg4b-bDhMbUfUfIb/bHdlfjfug<YRoHd6aSd?b0d-be39aui6aWj2a5asifeefdcOh4aHa+gA<a.jc6hWhx6bhahWhti<br6albkf:hNdpiC5FnBb@bGJ;adghfY1pbub|bXF>b*pPf01yg-avfruXf5hhc3h:gEaAe4g\\\\{hyhSf9a7btd-a5b.bB\\\\{yh3a=a9a7bJ0s3g53ecayh53kG3a33iha,b9a7bn[3hmaTiCaLh9a7bHYw3aoa8nnhvg9h-byh3ak3awaMi=ekfyh3asbzhEa3ajc?am5ctaLgzhCaRf6aXh>gOgMh:<@[W3Erag6atfNhVhwh<b3c-aX8a,8aia2h?aRf6a95e/a?h=h6a<bxfig4oKb2aauIbcpjf8fwbXcjc@aCcVc6a\\\\{?a&aub5c5aye=anbSgybrh5a\\\\{e6a7bJgHawbXR<bsa-b9a9b9aDeSg-a6a>ao3aea@a@aq3a%a@a0c|b9a0b9aH;7a6aH;Ia|b>d9bJa0b)3a#a-b9aDe9aUmJa9bSgnbJa6a|b5a,bHaD4aga/hZv-a5=a#aau/fau/f6a8b5a1btb*e-a=l*bpL-ay3aba7y3lka=l"));
$write("%s",("jd|e/bHdz4aua8b9a7b5aMaJayb>aSpU2??aAaHajgJadsU2Ja-b-a\\\\}c\\\\{c6a@a5L2b.e|bMd:aLhJaub5a-eMdL>4b-bJa3bjc?9ceaKh3ai=aQ7apfThRf;aYcWc=lm-,eKi;i3jok\\\\{ijjYj*c\\\\{jtkckDh0:,bT=tCX7gbW6GnCy8nE28n1s:\\\\}wbtzBn3*cm.b\\\\}EyB-Lbb9IO,Gt\\\\}/D+O,zbRt9A@mM=;p,btCC-xlSzgl>a.k=akmZxXXhb,W\\\\{@dbSz;J\\\\{4DLQI+kfb-lMtozlb*bY|Z<gRkbLm?rviLOJjJZcRAaMz,:/bmbdb\\\\}bDrjI=atbZ+y7nlmH;Lfpln?t7\\\\}V|iB:k@ouFtn;\\\\}Qp<a3NFaHw*v4bXaK9/bCaw0H7ttwo1sDY/bS8KzMdYap?Y:gARXH+kbVI<z:uvYbIAaXaSvWaGSRa5\\\\{xI>xBl=a1NKk=5-bXAmbv60bP+DaszhbDa+mmt\\\\{u8bwt.242\\\\{zOa1lRkzMWab7e;MH|b7\\\\}J7V|ZCPk.5-MJo2g7mylp4>aRXQtds1\\\\}TZenDq;<lpfbWaDY0NNJ8NGHEZ[T?Cba7T?Nda,43H5[H5Cca36I5Nia(ntnirpnW4Qba2rTOba)D7[2:[2:[H5[2:[*3s#emt.1Q9lpG/.?s-UC.b;@Rt=abbubm-P.NJSaD2\\\\{O+@eTa\\\\{Dahz8Q.bDrkp4pznWaew+bpC/bM:,L\\\\{bPk.ofpD/wt"));
$write("%s",("Pa|2|\\\\{<eTa3ESaYaz4b4Z+ul1*YwJ4El7l2bqmqYMEibEaRXzk<a?1k+Psj2f,od:2|Np4In/+ytjn1bzkfr5k5b42LycVEa5bM:a7U>om+2rrT@mn8rP@iCmnH/K@-?E6DaPa\\\\{|S\\\\{Ea>aVC<aftdbXa\\\\{1mn,bJ7DrDa@a8@b+EalSurEaMeYa\\\\{t/b,x+@\\\\}@u3>ak+l/PlpCG/WBPat@bA42YoSa8rPA/bS\\\\{h9m-G:.oWPDaTmDahzG:lbT?R?OI3-N?qEiB18yk2lEadu>a@xG?Dazl>a@xSzc3aNcG?Da;?MM2lEao:C5*GUaCLh,O,dbPaEahdfQubNlIE42h<\\\\{.lZSa7;hbegKQ2lomlbswwP;u;pH/c-g<lb*b2t?kLv0k8ngsjb7lZ>lb2bJ=lb<a*bO,.bOklbBk=v2lyk+mcmzbbqlbp/PaCa-bJ=+M7bmrilgsjb@>Da*rqHCaYaYr?aYaYr-b>MSzDl.b?qlbGtDajbD+cmGtDa6dY|ib\\\\}>dbG?cbdbG?:2Jd:p=am-WaXX\\\\}HxlE57b[k0bb|p;Om\\\\}BWz2bJ@|+,lbq2bhD.1crXl<a9bv|3\\\\{*kglS==aTahlZQz4Ya*kwvGsm|ubYb=aTa;nAaBFhbsE-kf+/IQa.1+s+nUz\\\\}=Uzxf1K?awmUz\\\\}=3l.1n00bD\\\\{<n3l?aDa0bLE*DwmhbR=f4U>m\\\\}=aTa<JUvsP=aTa<s<aZ\\\\}:-1l+s>aIqAe"));
$write("%s",("n=WbOahbcx01Q6EaIqJvp?2bD1ub\\\\{tFlBakbjxeb@aP2nf9<7<*bZa9wi9zb>8H/qX+nzFH0EacCZanX\\\\{tVaCaoJH8PlZ.vb1Xm-E-pZPlY\\\\{jbO@I>mPXa0bN4z3a7+kD0pCcCUaCaK44p|b<aAlG::s6\\\\{d+Dambz35=3WP/8DgIDa?aSlN1Z<<aTa1zib.kAuTn5sYaJT@pB8N93bstab98Moi/YaA2kCO@I>D+5p\\\\{u+b\\\\{b4|SB9HBn72>xQp=pHsSB9H9ysPbb0bRt8b>G3|h=ov=r\\\\}|BF2b7\\\\}v|ebh=4,k9Idab<w3bxlcb3|/bEa2Bkbhsc7lbo@*odb4s8DIO9mA8R|eHD9I6RaEkb@/TQ@G+uv4NZlCaBa5btbwnLoD91KGa.clDvxNmB2QkOk=s.LW.rB84*BL|hb3bLnm\\\\}W*s7hE/Cu,Qa\\\\}@z>v|71Y:jRP/UCOahfZ+*xD/cNYa;X+rtbYa:uP0tQF3hfXaWvK.=a\\\\}b4bGw|GP/XwK,+A4+S\\\\{Wn=?RmpG3/JL*H.UX-\\\\{zJ\\\\{018-gbeb,uW1|bZo\\\\}bVwP00bjbASlhyboOsUFzDrxt\\\\{mxAP0cRz16IZ1??Dt?tJoVaD/+yPt4bRaN-ebabC53>ubBFvxWS0b*b\\\\{1BfbIgugUw4Zagr>*oOwUe*c7oFLMkb|brlRam-9ur5z-EBbBQ6QrebKiPGIOPa8QYcpCjNNaX<4\\\\}|c?0lbv<wWyb?0d|3"));
$write("%s",("d,b<HzbdC?a8:FzTrW-EtB.,b<H@oA--L1n7R<HBtnW#3awgUag|8tAnoCd=cblvgBmOPvQ6B4.2Yrib54Oakbf1vbYe\\\\{wzbzb<sF4cbQO2kzMgsC?p;gqH6X2pwMsTaKlEaY7x/H7wwOlQ<dbPD0\\\\{gb8w6wN13w314xKyY,314x5T66qZC|KGyv\\\\{hrTe3dp,b?aVK1q;Qzbbbgb+/>5-U6>grdg*bRa@wEQU7|ozoF3mbJqZzgn74jDel/nxfAa2PiBc7.bTmm+/oa:>HZacgkP\\\\{biCuJ.bCn0s.tVayvuu,b1t9BPaI+tz2b6/+7<aCnvbF4GOiCEv;rPt8m4lys?tIncMiEhjWv3;mb;r2RDvGKKN=a6PP.58k/O|W/K0\\\\{+J,+/uPa.QTNaeb,sSamit\\\\}D>8bN</llqpu:n..<zpuubl.YM2tg2gb->AaxnkbqZx;bthsb==:3Fpwx7y83b\\\\}@2\\\\}GTUaul3L7lbI=adE1\\\\}y|vb.oq39nq,.q<1AaLw@DPyTpYsIEa4>2PyQQr3K/-bDv,jDq7bw5Ra\\\\}/Gl=aQ5iXlbkp@kuy2/PrOa58\\\\}b;J6.wP?n\\\\}/Gl=4wxu3cPg?u/bavOa2/?24txfiI5yA3xtZ/I,z+.b>DwP-,=pFawpA\\\\}31w*Y7avP2zMT*@aNaEatwPaUvgzvk0Pibd7P.Efo<*k1s?D?ZBn2omO-ncbB@4bNrg8B.HVOYGmi\\\\{B2ybc31@tbQa:\\\\}"));
$write("%s",("//Kq:8N6iy+rL80qt|Xa<k7h|p-\"\"),\"& VbLf &\"(\"\"U;Z\\\\{sxf-7ybFaa1qupIa|=lKODQp/RxOm<BjCXX3>n9?Dw8-ZOa=nawfb\\\\{bxbksNf\\\\}nVTFay2V?j5hYdl5HWB1,.\\\\}gIVTGXtm3M\\\\{bL,=r<\\\\{QV-7DEng\\\\{bub?=HupIkbzbb.F|Hp4N@9*r/n+r8y-mBB?1zw5b\\\\}bIQfE>aEI,zHqNx9b.F|y=9Bphsxb98D/CvabXAIm9/6bOa;X3t1b+bwbiC5bJt=3Rv\\\\}br|,qY0f-pIKl@BstEekO9.,djDRa=32sNU?a5pPk1b*bSa|\\\\{n/=qUKYD:q\\\\{zcVz-qoLyA:4rpum--n<rPa2b72Wv|nL1asFayb<rk6>>1XH/Ra5HPa1X,baJ\\\\}bg@LmVp3GY\\\\}1uPat:F\\\\{xbcRi9LiXa-b0ofQhrH2wb0<bbm:k:Oa6\\\\{Y<\\\\{\\\\{y\\\\{w\\\\{1rkb4b*y12nKa\\\\{q3krkbj*9,TQba0+TNZ0\\\\}+b?az6cvQH.bClq3s:8M>Dfp2W;r2bw4ln>tGabQ<npI?aO\\\\{H8+b8bhbW0n9u2I99sc.>OvrRp.>6F+b8mGynu/biML19=HU\\\\}M4As?/bfpYa4AUa\\\\}+\\\\{bTmjDTa05|ni9?*:pYqoWJL/bibY:MrgBxfm-SE\\\\{b?a85Bab5WDRn4N:>4bRp7bOJe+xbBal,w4YkH87lRa4x/6szguiq/kn.ybqzbbm?=5\\\\}"));
$write("%s",("5bbyb@M->wt+BCwAzL58-*rAr8mhfC5A5WS5d|oKqs?q:Hh2gZa9k1pI8RCu<t:LeI5rxbb6qBa9/;\\\\}Nr5q7dv?/8af.rdC\\\\}5c:0zmr>>ApKl+ABa;I*b3sLqJq/nkst2.?O@.b\\\\}4Naa|dq:Jqra|A,LvXk@UApVxctxm28HJfbunPKHzZaqd=5Dh3bFnG+<6*2Fnm-p;c7p;w;\\\\{btFxb|bEP-b,q9bUazqvozokftCjbY-kbV.zbdb.myu/by7f@>5hb@zyQ7GVaP.1DVaf67bu3cbCKMpHu?0EI\\\\{Rwb0/owqMbq*bLuww,bfQjnS7Q*I<Vb5NAKd*1bk9m*B903mnCert/bPDEBnTR??aGa,//oE<rhabZ8qERm7dEpjbb5F2<e/bVaPaPs0PdgjbLnsz<HC|ln.y\\\\{wE6FaN4gbwwgbEaPm@Cyb.bpw?uszFaG-6w6=VEY:;Q<zYm3LI<ubysc+vIuumzAambfxYx7/m-jbtFd|GH3/nn?6EaPaVadOxo3xG+H||/jb>/\\\\}bqvxODa|b|;bbPRf6k1VtWKEewFiBuPfGI5L/wbEPy528e*Vkjrx.c,nh.R2RNa*/|b4k4b\\\\{n=aW?CK/bG\\\\}eIVaf+Osf+vrRaFa|?;I\\\\{p7mL/I/K=@sEa=pG\\\\}z/Ga4v,b<nSqe*B<Ca7mF4Ua@aw|S.A\\\\}:+Dq*oB1IoQlWaAa|t4p4*V|T/q19betRx4-Hkp<8:iyGmfbLd<nkCcbB9WQ"));
$write("%s",("CatbSaNaZafbGmy,|beb<2t?Teebsz\\\\}b@a*1//.baukBj>3b\\\\{2wto9q6Uhwtj6-bu2mHbb\\\\{t|?>zlotb,lzb;qv:jQVISq@aAawQOa?a9oVf@a|>IuA-5bc*g@y0<aY6f.-yBaSacbs8v-izNa0tYj54WqDzOx0nGaDIdg>i9umbG=W?3by2Y1DrqvDv|?vnlnqFuFmbGmFJdP:+@+LwAaOa0P\\\\}0.s:qQaWaWaEe2;<+AaK+RaAavD@\\\\}8<l<i/KvAKPaL,M\\\\{57kbU6Qa6=\\\\{b2lf\\\\{hbG7.b>a:,jbu2<a18W\\\\{PaNmWaOaPudObOK,Na=N;rV5eI*x0\\\\}=ad+M+\\\\{bJjcz@wjBTa:wYM=N1b6;A28:Iy:ojCebQqvn0BP\\\\{8b+:G2xbgbhF:s;qf-Qq1bFJa6Z\\\\{KqcmOacbNavbDqebkn8<;3W0zbmb9s;s-bdbkbtCFa<avb+,VvP0QaSa.b6lSaGae-x7P<AoZ\\\\}-uq4UaHnz-e*r\\\\}Eaar>a|b1x-771XaqMdCPH6+X41r,ePqRa/b;\\\\{xu-rEaMHettb>aiba7jbWa+rEBbbdb?COabbYa+bLoCl-q1kI7Xahd3dvbG*Qu3bbbfbCnFaNaYj.b9bAr*n\\\\{EYa9/0b=t\\\\{bPKKfstm?y|6dF\\\\{28MkCt*1mb6bebiqm-nuFz;J9|1bTaZ\\\\{10RaC42b9b|b47FaUa1v<Bim?C\\\\{n\\\\{bhb-8Lo*vzqCa@s6bl"));
$write("%s",("b0baJf,cb9.QaDa<z5bcM2LK?,bUnC>Ap-mh7B*-e>a6-MvKzjxIEebq\\\\{qvNrzq<L:L\\\\}b8LE2>D|bBpYpw44f3t..fpQaeb0sXwabjbEa-b;J-b6b/pFpyqf7kben?.NJjbAl<aeb3bQqNfbqzbDaCagb6rDa9/ElB1:KZa|bvmMriI;zolNaBbbbRahqB9wK-KubA.M/bbfrI+42*5D+z7xn7b=KQa3beb6+Ar9KXufbm-=xXeco\\\\}b1nEamn@aGh2;,efbqvvb2K6+.?VahKmbubKwmb*Kv/qvxk2ky0Va@?+bvKv/wqrKRaRlqK\\\\{bz\\\\{wKvrg07b>\\\\}|f7bkyMmI9A.zb2k.xA8B<HlBad1tbtuhbibZaFp2;j2DaPrzb@669I|>aaJrF1bXatnTqWqew46.bPa+b9\\\\{\\\\}nC0bb+A+zx\\\\}>>-bhb?a8bkbEazbM6H/I8:\\\\}>b*1os2k@amtagymlpt0hzyb7dd>zb0bGmRaB9??hJBaV5Paxf\\\\{zUqiq<amzmp4qt\\\\}>52bNaPafbNn08Ag9\\\\}kb<1gb*DXxvbv\\\\{ib\\\\}<<90bTsNay?K4I4FaxfjbJ=Va.qRa+E|bs,,bBaWk/rhb?hUaTl<a\\\\{IwbT|Datbl1lbDrL\\\\{180y\\\\}8-bgsxm8bomibT96bNrI94\\\\{<ajnpFKznAH72b<a|?*b6/YaGGGa2Hy-zbgrjb/b<@?\\\\{eb3nbg/b1b=ahBbbfB5y//rs=+VaP+"));
$write("%s",("9iyAGwk7@D0+9=Oa9\\\\{tbrFj2gbYa>ajn4b>2xfebLkC7P,exZa\\\\{bI|hbCaMs<B01Qa:vwuXaq3Cw8nq<ibDh*yz6>aJ7c,Uy=1:1M\\\\{/b4bx7s3q34|Caa?ds>8m-H/MxR@1q\\\\}pzbrr1kcgpocg4xNfW.XwP0ZaNkQ.XcW.jqR|1b-bjD-mUa0bWamb1\\\\}woxbCaM\\\\{W35bpsLC\\\\{pXvebEa0:tbctOyv<s,PaYaQ599U;F.-ktbv<E2=@XFz-NFAaFFJF>aYqMFXaKFc*pvr|1byb6jt@YaNrMpqyz-9b2bEa,qx/DFwz>D-qB=5AN-2Babo,<pfBnnNlRp>8==uo69af/b|b8b7\\\\}|n,tu;sqjb=a-E6btbU3ebH4/bYa|v8b|bUa.b1\\\\{hbc7Faxyebj2B9wb.,Dh+b0nm-GvybbbqoknApFahbSrQa,<XaK6SaibDtL.5.mbtlR+xnwbH8*bIor3QaD*S0z+|Eyt.2ZxxbvgPDHfFr62\\\\}:Q<Zp\\\\{blbct-eZpm>+kN1QamEGa\\\\{l1Dwl4b5nzbNaL,-8?aB6Ca0t1DZ\\\\{V|y\\\\{@v8bVaDa4*8b/uXa6pvbRDPD3bib,bMDltJD|/1kYaFa=D0</*2bN47btmGy6b|bV1<p+;3<bpEaGar@ibV>H+6rnCUao2uDP0Ea\\\\{bpyUa0-Qr6-n*N?|*=aXbpplh0:mb-q4f@a2k\\\\{<XlRl?pEph=0r?qm-5b@avrR|:\\\\}lnjb9"));
$write("%s",(">1wkb|d8b=@qyW.XaxbO06t\\\\{bN=I>I.a|rm0zmb\\\\{b?oc-zbxf>Ccx>str<?Qa+b+,|/wnrlDoI59m.;|0fb\\\\{,d|Vvyscbtw1r+q=aFlJo9.mbbq=oQaV9DuOqPaub>xgbAkTa..Ra>>0bvbTaFaOa9bClPaFadbDa\\\\{b2b>@Q:>aR\\\\{I7pBubOoz8Yb\\\\{byjl.\\\\{bOzRsgb1siBxbxbibK=:dRxzbCl7d?rxb/2dx>awtd6vbGt\\\\{zInYa\\\\}bSa*wRa<aHm\\\\}b.bubOa:n8nvbU3<vyyL1Hmlo\\\\{bv:?0*w2nUa=lbzO5mb2/0qQa|l?tOlybVaaw0q-bab07:\\\\}2pTaOAjbZaQ.,bIq*:>@XaCnqrCl\\\\{f<aMstmZaX:yjEe>@Va|bYaQt*pfbenvs1bhbI3Q9IrI<gu-8oi|y2b*bX:o<-6IrQa:uxfK4/rgrilx\\\\{b*C4RaVa|yDvgbhfYct0Oa2bnzb5G1<elbAnu.>@R+?\\\\{xtctM@xf.b.bTaLuPnZ\\\\{\\\\{ddbHhsdxb@acxf@gb\\\\}bwsslr-kb-bAa0bOs3bVal/Yv9>,rV,vmdb-bZozxuoy\\\\{wb1babGhDaWaVx\\\\{.|uwmzbhbYq2bdw\\\\{qzbOkPaV7xbWab\\\\}cxcbV9Gat8Tmvbol8-hbabTacbbig+kb>aub+oox5bvbpqmb<>ow3?mbCtmb<?vbMyfb!![2aba!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"g3b[2lha\\\\})1(f\\\\{#*3&ga(f;)0,W3MZ0=akb5>Dr4b2g\\\\}12?PaG*/?h,\\\\}1+b3b9p>5,bdb|bP0lbwmybNa;rVaBaU>osR6Y\\\\{-bxfg?vdlbW\\\\{cbOaR>M9wnPnW/Zx1khfI5od7llbyz9pJ=R\\\\{RaBaspubV,6bUa<aablr,bg0a2gphf9podL\\\\{dbI2;<F45bw\\\\}xf28tbbq5bwb4|+wYaCt7-kb+wHsA0bq\\\\}ocb9pB<.\\\\{i7fbu/dbfbebcxn.Mt.hDrOqvsIokvxb@ryvm-0bo-7bEaxyFaTa4dN<xl5pmzyu6b2p=a1bO=Ea9bcb*b3b=5Gar1bbZa96YaA3YwA.ab8b:y.,+beplzDau;*/Ba-ytleb-bStcw\\\\{xV<\\\\}=V<xfm\\\\}?j\\\\{zU<\\\\}ba8z\\\\{n9tb:ykbs|?jebgs0b*pK\\\\{ub6b2zm\\\\}St0vm0eb63PaoixbBl3bAt,b\\\\}\\\\{3b8b+bEaM4ebb/mbUawbWa9i,\\\\{G*bnXaZm/<HtQafbEa3b|bNpkn,<Mswb3bGtI7@amb1whzQaxfGuBk9bvb-fK9Da1bEh=aE6ibq6V,vpPatbu32b:88btbUa-bBazx5bWkPmM\\\\{-bebxf"));
$write("%s",("..WaAkm-R\\\\{lm2bA+H\\\\}2bz\\\\{/*EtRlH7lb9bLl1kksFl4;jm>amb\\\\}bwb9lY51v*/o-Y6BaruI2oohnMzDkPa,bxh|bSa=a4k/n\\\\{16b3begwbybzb,b6bSa+bGaRc0l3b1\\\\}Ya7mvb,bQ*<aEaC/-7q:|:\\\\{8VnjbTa<k:k8k6k,bPa|bTakftmgobnbb*bQv27U.,b/rvob\\\\}EtPnvb.l6bX8>ar8>aEaMzStDa94|gkbYpybH\\\\}-+wdc:A25qC\\\\}bbL,o-ib7b=x?aybc:Bfxf=agbwbAag2/bOa>a1bl8UaR3?abbHkv*9t?qa*CeV,Zaub0*Ba+vU9m-B.ibibXaPaMd4bZk<aDa+bZ\\\\}7bE2tbPa\\\\{b<\\\\}*b,bmo7bU\\\\}BalwEaCaHmG*2-M-o5c*4b+xTvhdvn.ba\\\\};kTvnu9bJ7RsA3:-|v\\\\{x;\\\\{0bi9=pwutbnq-b06ebzb7bewB4/bPa3blb05vx,q|-Br4uZm8b:sub96@aebhbwb6wyuOmBp,uZ0Oa=a7bhbubV+Ysgb\\\\}0o.-7cbVshzWaM\\\\{IvBtTa=ad16\\\\}0bUa\\\\{b7blbBaPy=azbZaOqTnefVaNvb\\\\}xb7b-yxf<e*w5eCaL-b+*bFxa5n*ub1rVu8yw,wbhshq*e/z5fnyD*WaXa1rm-bbXazbjyM7K7I7MokbWa@xibjbjbkbE65bPacb0bLvibN6GaQ0*v500nJ-?.sv3-Va5bhb|byq/b4"));
$write("%s",("*hb@a0tyb*bv*+oWx9\\\\{Ba0b.q,qhxw0ibE,Ju1v/*D/a5P.2bcvfbcbj2bb/6+rxb?twb?lab-6db3l2b5.Pvlb,bv-L-cba+il2babzbPa+s,bjb*eL,H+VpgbTadbM\\\\{xb>aiz=ak,A\\\\{gbT|BaNs5yTqyb\\\\{b\\\\}r5b4-=vxyov1oZkjbHuOqW|+b4bR,mpnp0btb:w2,rsMtBtCnybhbenmb2btrXklu5b0sCat2dlibqoGw+bClcbm-Ea0l6dvn-t>1Xq2sdrimww,-xf*b>kRnTaYaQaf/dlr|HlH+FrU3G+ub>epdPy|bcbwbVaBvepgr2g=tMpVsWaY3ebyqVsV|c\\\\{8bktL\\\\{J\\\\{1b/14b|32b>-<-yjkf|c:rGa7r?a**,b@am|@pxffpdp;.j4R3jq\\\\}b5bznmbebtbtbMl1bbbhbZavbk.Mzy-GqcbGhb48/WawbGtTaxfS1lb\\\\}bdbr3xyTaRqAaqv=s/bfbDa\\\\}b+,r*Aa7.Srm3N\\\\}L|ab\\\\{b,-9lQx.o+nVaTlA\\\\}\\\\}bhbSc,yabYaZaxbebFaWahbzbvbsm4bBvV1o*pv\\\\{hm-6gvg*bStlb-bElrxRsvb7bY0.\\\\}cb5bRqTa,-Wqbv\\\\{bStvpYa0bKrTm6bXmPnbb,-F-lbGaPw\\\\{bXa6\\\\{|-4bF.DaQk1|cb/babVpNaqyfbIp?-=-+reb4bybdb.q**EekhFa0bEa9o1cwb4*Rk6\\\\{Oaib\\\\{b6d"));
$write("%s",("Mlgb<nQa*bhbe*SaBaYsVa>alu*b8bDz+bdbdbOaEl-bNa?.-b\\\\{qitNa?p*10bLern6b,bQk@akbBnVa4xOv6bjb3b@a2,i,sz4b/,Ru+nZ\\\\{ZaYqX|-b0b7u\\\\{dAuI|Gavufbab*bWaO|q\\\\}/bFaX|2,<eOaNacbA0\\\\{b,whb-bN.O,|b>0.bZzdbybGaE*m-ebqn4b-ntbTaXrIp*bUewb|bCaDa;ry-kbNahzQqFafbXo1*rhm0*kFu-yUa/ba|zqQ*Rl6\\\\}+bHkebub5\\\\{dbZn<aQa0rRabb5bWm\\\\}bYu/s0b4bctkb9bwbubDa*.ubxbkbdbr\\\\}Utu.hbgbW*ubXbWaGs@aQaUtUacgXeTajytbLk/kGydbwlUac\\\\{Hf=aTpzw+b\\\\}b5x8yabGa*t*qwb7b9bDa8k=nWr+bXan.tprpqo6gBaD/\\\\{t7kWaKw\\\\}bVaIm;,ab5brpzbo-V,>thbPa<albLoWa2vg.Fa,b>s,qFaZav/4bxoOl-f=pVx2\\\\}mz5b?jVajb9bfuwbYa.s3b<am-xfWa8bEalbgb?aMpQ.abiqSa|bmze.ZmLk>aFn>kSaVambgzYambLo=aMp|yYcKu,ztbNnkbFaTpdb4blv=s8b=axb\\\\}bPmAaabyb6bvbEe|bO,wx3|bb7bKrDa4|w-cp/bwb6bZo@uybtb6,zb,w@a=aFa+bY*rtCacm=*VaTaiy@sabbdy-Ragb/pP|Tlo-RambTa<a|bqoy"));
$write("%s",("\\\\{Tv>amvmb1bmb4b0b7bibUakqApW|?hgu2\\\\}0\\\\}zb8bbbM\\\\{zblpZa9b8bZa6g*k*bAad|vbIxdbAaQakmuyAaArAaNaRa?tWa0bO\\\\{3d3b*xWlYxjb*y:,Lz*bybwbwbVnZaUadp|bRatbAoYolb>lO*=aCe6,dbm\\\\}UvxfDaV|6bcbabAalb2wWkvb|metRsr\\\\{EaZalbmxy\\\\{Oa4bkbabH+gbj|qvArmv|bibHlUaylafybQaFaSqBay,@aOmKy?aOazb@a-bfb|b<zDaJuQ*\\\\{b@a5eYapvzbFatbCkBa\\\\}vEe4bmbzbGnBojb+bVa,b\\\\}bkbAxWt>a6fSrFaBgdbPrFa1zgnGh.bf+*bBaw\\\\}RaOaWap+7bvbjbmt.bUa6jQlXambc+8bWagzWaSam\\\\{;mgzRaab\\\\}bxfroZaVa8bRsSa\\\\}+Vs<v/bSaQaEaAaVanqOlm+0\\\\}EaabQl@aMp2kmbg+=aYeAsOsWaPaWa@aSaEaib5b5b,|Ta2oAxAacbY|9bvi7|\\\\}bfsItabJuC|1\\\\{TajvYatb,dQa7\\\\}kte*|b6bNabb-b*vdqnhm\\\\}vlZajbT|8b8b7ba*i*-fyo1b?nwbAgwocbk\\\\}Oaabh\\\\{Y|jt\\\\{bwbYy5b1bYa6qo\\\\{8bebBa+b1\\\\{jb;\\\\}8bXa>aab>aVa1znh9bgb=pPomb<ayb\\\\}b1y=a<aGm\\\\}bibVa3|zw?p|xCaVacbxb/bImSa1bPakb"));
$write("%s",("yqtbhb\\\\}b/b1gwb.bVaqmBaY\\\\{Mmr\\\\}-x+xDnZz@|*b@aUa?a<awbLd|bNawoudtlibfbtbGywbudEq,q3|,x?a3bksAaYaBaibTa7bcb5lAa/btbVaxbmbgbib@rwbCa2lybns,bmbZzDaRa,|*|Sa<aRatncbJj?wDaw|tbabFltbUpFuRakb/b*bPoOawbTa4pQaQuabgbqigb-b+bfrXa?awb/bszib6bPaPrlbQshzPaPa-bFawbNa<aFazn9tRaPa>a=pOa7bktFa2bCaUaExjyUadb,xmvlh-bWa6bZaZaal=q8b?p4bruab|bjb*b7bbb4bUaBlAaxbyb2sUaablbxocbkbAaozubXakp?a\\\\}bub;rebVaSah!![2aba!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"g3b[2lha\\\\})1(f\\\\{#*3&ga(f;)0,W3MZ0j\\\\}b\\\\}bbb/b+znmUaDa5bTabbxb\\\\{b+bhbhb*b-eAa.uCanz6bamDaibxf\\\\}rfbxbPa.b0oOa/smzybvbub\\\\}bwp2bFa*r3rzb*bdbrzyz8bFakbjbyb@a+eUaFact?psz8bqzfb0bBact8cUaNauujbBnDakbgb0bHd:pmblbVaVaOa"));
$write("%s",("@w5oauDjXaYaWa,bnsybAavb5y@scbXa2uNa7bWars3bftEa1y/y-y+y\\\\}yJuHuFu0b5xxfxlJubb3bup,xSazb8qykAaebjlmbxfibSaXaRa8bwvZhAa9b6bRa|bRtAuwo5b/b|l5biblbYacbbb>eZvnn.pExOoIlhb>a3bXa=aSaWaHoOa.bXa+bDao\"\"),\"& VbLf &\"(\"\"u6b@bkb\\\\}b6bDvdb+n|buuRattNadbfpBaebvx0btxebbbWa>nkbQa\\\\}bGvebqwowRa0bcbStXacmXaZr\\\\{bPaQo4b*bew2b+bkb>vHnub-b0s.stwUaUaib?azb\\\\}blbUa|bHvHuXa4b8t1b9nRweb1bxf\\\\}bvbqu.bSaCaxw0b?acb,w=s1sBa:v4aFjZtib\\\\{u7bvrFaEa=awbPazbwtfb6b2bCmsoCa2dibubxfTuDvtbAaMsQa,bewRv>aeb6b+nkb7bVa*k3bSa\\\\{uxfafGuwvdbNalb9kubtb@alb\\\\{b*bXacb2b7bZk8b6b-b>aQa>akb4f6bDa.bZaQaCa1b0bmbSnQa=aEacb\\\\{bib1bYkhbxfabasjb-b8bwsZaAaMpmbBawbUa.tUhFaUk0b<oyb?qkbepbbjb7bPk=a3bNaxf6gjbBl8u.iwb?aXaOaMp3bUaYclbvb9bGaopmb9bDnhbdslb8bAa,babmbEaVp<aubQkibzb?a4b9b,bXa3b5bCa9bXalb=a5qDa\\\\}kAa-b\\\\}bmb"));
$write("%s",("WamsRtmiubgbzb=adbxf8b\\\\{bVavb?adb?atb0bsdZaxf1btppdZatbslDawb4a6oyr+o*kuoCa=a:nYagb|b\\\\{bYa?aPa9b0phbnqzbkbdlgb*b2bYaNa*evbXakbUnCs|b,bNanmCatn.b-bZaybcbtr*b\\\\{bybxfFa>rvb*b+b,bOaCakbMo|ndbebjbAaBaBp2bbbbbNaab6bFpcbzblmxfQawsulzbpd.pUa@plbDh>aBpmb@aFabbXr6bybYaubab+b5bybXa+mBalb1kubPa1b7bBabb;pFahsEa1bZa-b3b0b@aVaeb+b<a-bCa\\\\{oAaDkgbOqababcbYnybRa>a4b<a=a5bYafbgkJqwbSatrBkFa:q=aCadb=a\\\\{bzb5bFbybgbvbUa4bZambwb|g\\\\}bGmPa1qCaxfNnjbBa|blbjbOa/bDaUaEaxbAlxf|bab7k5bZa*n|b/bkbeb.btbjbabRa\\\\}b-b=l4oZa7b.bBaFa|g,bZa6b.b\\\\{mBb?a9btbVqcb7bNaKd7b<aafebgmxfwb\\\\{b/bdb7bZa0bXa\\\\}b+bYa|o\\\\{b1bdbmb+b=aBpVatbQp1gdb>hebQa\\\\{blnlb5bCjcb6bwbXa2b6bWabb\\\\{b.bOaXaabxbAajbGa@g\\\\{bmbqqbb1baqdo*b:kubkbIn5b|b4bdbbbzbabPadbeglbkbfb,b0beb\\\\}b7lgbubAa>afbwb4p\\\\}b3bubSnBaod\\\\}btb@p,b."));
$write("%s",("bmbzn|b7b0bZaab0b-bSaPa4bEa4b8b/b0b/p7bXa@aubTalbYm2b,bQaxbNaVaVohfvbmbOa\\\\{bdbYa7bxfcbjpubcb\\\\}bOalbxf\\\\{bWatbyb3bOaAaFa1bWail?a\\\\{bpo4b3bcbgb,bjlab4bLn5bRa@a6bFa+o4bxfyblbTagb>bNmRajb,bGa7nvitiHj=lvn4b+bTaZaib9bibWafbbb6b4b,bWaCaebib4bSnTa\\\\{bkbxbRavmFa>aWaznxnvnPasnqnonSa\\\\{bYmWa>a+b*bPa0babQaUa3bDa7bmbmbXafbmb0b0bGa\\\\}dXaUaOa,bvbClRa,bTaNa5b3b,bxfxnub8bib-bbb?ambSa\\\\{mxbTa1bFa.bWaFaebXaQa1bfbFa8b2k.bAa8bCalbSa5bkbYa8bDa9b-bOa*bFaQapdkb5bOa1bCaAaSayb8b9bzbjbRazb2blb/bebwb2b1kZl@bQa9bfb-b7bSaab>h7b,m>aNa+btmUajmhmnmlmVa.b7bPaymTa-b7k0bPabb2bjbNa3b.bkbRavbdbhmvb<a6bBavb@aYaEa?a5b-kcblbDaFaVaAecbhb6bEaDazbWaTajbUa,b2b?aNa>aTafbibOaYajbcbib>a/b\\\\}b4a;lGjIjudxfEatbDa/bhbNaBaDagbfb>aYavbRkPkNkxf4bDaYadbzbXaBaabwb*bCakhZaFagbVa6bTaQahb<aYa3bwbwkXk?aQa6b*bkb,b"));
$write("%s",("ibvbVa0b.b,bebYawbvbRa7b|bhbRaCa/bjbhb,b*blbhbTaxbzbEaubyb7bdbCaEaybLeQa4bSa>aDa*bibBadb9b*b-bEa7b6bAaEa<ihk|jekNjpjfjxijjaj:j;avjbj?aZivj\\\\}j:j-b<iujCa:jwb\\\\}c<i4j8iOjEa-i*jTi:jOi4auiEj9aviSfsi/b-b4b-a8gubofvj-jqj2j,i9aEaOavj/i-iojue:a-bjj=aAapjsj.ipj6iej@a<aydViijgjjj@i-a>iYihj:aCa8acj>aAa7i<iBc3iIiAaAe7iQiliyiBi:iBa*c=iEi*bLdqg,e5bxb*i;i9i7iyi5iOa*i1iBcAa*c\\\\{b+i2i0iFa@a-a,i*i|i9ayi\\\\}ixb8aCa@a*c*e8axiHa8arb8a8a2b4a4a3aRf4aNd3bWb6bfdzbxbubjcLfMfKf5a,d-a\\\\{d1bGb1b7hhhAh;g?a=a0hIgefhcXg=gVg>aBaKg|b|bvbag.b3bzetfWgMgBa?a3aHbXb8grbIg?a>fghCdehDaAeKg2b3bNf,gid:d-aue-b3aAaCa3aKa\\\\{b;aqdwbhfIa3b1b2g,b|b0aefbePgWdNgDeKg.b,fefCdWfUfSf@aKgybIgtf<fXd<gBaRf5a3b9f1aCd1adcHcubwbxf,btfVfzfTf@a3a1bhfwb+b-aYbhd/b8bifXc;a:b6a5a-b;dZapghd5btgEf3bye7d5dNf-awb-f3b|d;a<b:b3"));
$write("%s",("b-a8b5d,bxb2b2btb;aefWd=fPa;f3a>a3alc-aLf/b3b4b.bHa8byb2bpdtbyexb5b+bAbefXdyf\\\\{fce9cteHa6f5eGawfxb-b6d4a-a.b\\\\{bndMaja-bPaBabesfGa+b,e?adfGa5a5a4d2bzb;azb-bWb3b2b5c?a?ace-aRaYaOaVafbVaibNa=ace?a;a>a-aVaNaUaievbpbEaed7b@aCaCa?a>anb,eubFbzbzeMa?dke<bFaFa9a>a:b;aocGd+b+btb\\\\{bvb3b:dJa2b-abdocZbXbVb;aie6azcdecejegeoc/abeRbZd6a/aXdbeXdIcUdRbWdCdBd9a2b5aMdKdIdGdxbvbtb+b/bxb1b5a1a/aCdhcockc/aFc:aIaXbtb,b:avb|b+bub4bcb-bqdodmdHaebdbJaGaxb,btb-b8a1bxbwbtbxbUa?b|b3bvbxbfbocnb5aXb.b+cXb-avb*c|c6awb-bxb6apbCc7bGa7bnbIcyc*b*bIcwc/adcgcRbccac>a8a?a2a6a\\\\}bKaKa6avb5aYbVa5aJa7bHa=aGa>a:aGaCaJa\\\\}b-a1b.bybjcoc|boc7aEaqboc2bsbsb/ahcbc5anbHa6aRbdcsb*bRbobQbNaHa3b-b|b1b/bJaNa/aob5a/a5a9a4a2b2a4a5azb.b+b;axb+b.b2b-b.bvb!![2aba!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"g3b[2lha\\\\})1(f\\\\{#*3&ga(f;)0,W3M*3Hba3\\\\}4Qfa(f;)7E5Nda,43H5[H5Cea318368[*:[\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'4[N4.ca52E6[E6[\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'4[E6[Q4[E6[*3[E6[E6[\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'4[E6;da901Q4Nga=s,y=zX3I@G[@G[H5[H55ea11724:[(<[\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'4[o@[*3[E6[*3[E6[E6[\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'4[E6[Q4[E6[*3[KDlca91bB[KD[9G[9G[H5[H5rda616xMO\\\\}<[\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'4[h@[Q4[E6[*3[E6[Q4[E6[E6[*4[E6[*3[N4xda292E6Oza=y,]99999[gnirtS wen=][c n3aea\\\\{)v]y3b&a(niam diov citats cilbup\\\\{RQ ssalc?E[-H[-H[H5[-H#ca44|;[p=[\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'4[V@[*3[E6[*3[E6[E6[\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'4[E69ba9O4Nfa cdln?8Sba7?8[?8[\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'4[N4/ba1D6P/a;maertStnirP/oi/avajL tuo/metsyS/gnal/avajwJbdategu9Rda104u9"));
$write("%s",("[u9[\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'4[U>1ba6P4Noa2 kcats timil.e?Sca11J8[J8[\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'4[5<0ba8FDOga]; V);iVaL>ecaL[uVapVhha dohtemt9Sea2972$7[t9[\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'4[N4.ea4031Q4NzEnga repusW8Sda494W8[W8[\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'4[B<0ca06W8OcaRQK>cgassalc.f4Hba3X5Uba7U5Nda,43H5[HJEba11<[1<[\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'4[N40ca091<Ooa(=:s;0=:c=:i;):HajaerudecorpP9[><[><[H5[qF#ca88S8O><[\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'4[N4;ba3pFPqa(tnirp.biL.oken\\\\{@<bianoitcnuf)Rida\\\\{RQ;Fam:[V<[V<[H5[p9#ca20q9PlartStup=niamT5[B8[B8[H5[H5~da115S>TM5[;8[;8[H5[ZQ#ba5YQOra(egnar=:n,i rof;)X5[F8[F8[H5[F8[*3t3a<0Z0Z/512152353/2/2166263=4/3141625>>914151:1/z6[h9[h9[H5[h9[0Dvea+)6,E>[<8[<8[H5[<8[*3uea1312y>[;8[;8[H5[;8[y>xka(taepeR.S+#>[B8[B8[H5[B8[#>vfa41310M5[;8[;8[H5[;8[#>v9a=:s\\\\{)(niam cnuf;\\\\}r nruter;\\\\}\\\\})84-)n(tni,]"));
$write("%s",("1+2%%i:2%%i[&6[p9[p9[H5[H5~n9ON4Qba0N4[N4Dba3S<PcawW19[\\\\{<[\\\\{<[H5[0B[0BvNMbja=+r\\\\{esle\\\\}Y5[G8[G8[H5[G8[*3tbavH5[68[68[H5[68[*3t~a=+r\\\\{84<n fi\\\\{s egnar=:n,i rof;i6[R8[R8[H5[R8[*3[G5[58[H5[58[->2ka:r\\\\{gnirts)f3aea s(t,Yaba)h6[Q8[Q8[H5[Q8[*3tbasG8aN5[<8[<8[H5[<8[*3tbaSBI[78[78[H5[78[*3udatmfJ5[88[88[H5[88[*3tvaF(tropmi;niam egakcapa6[J8[J8[H5[H5#ca21J5Nga(tnirpfD[<8[<8[H5[<8[*3uba-H5[68[68[H5[68[=Iuhanirp teUT[>8[>8[H5[H5#ca36RCOfantnir4I[;8[;8[H5[H5#ca13;8O#a,s(llAetirW;)(resUtxeTtuptuO=:5>[T8[T8[H5[zU$tDUL5[:8[:8[H5[:8[*3sdaS C88[88[88[H5[H5[*3sca&(G5[G5[58[H5[o>[*3sba KC[;8[;8[H5[;8[KC[J5[88[88[H5[W38iaRQ margox>[P5[>8[H5[H5[w>whaD : ; R~>[P5[>8[H5[H5[*3tba\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'58[G5[58[H5[H5[*3sqa. EPYT B C : ; AD8[V5[D8[H5[H5[\\\\{>tka)*,*(ETIRW?8[Q5[?8"));
$write("%s",("[H5[H5[)>uhaA B : ;=8[O5[=8[H5[H5[*3sba [2cN5[N5[<8[H5[H5[\\\\{>vba:98[K5[W38E5[E5[E5[E5[E5[*3[E5[W3LhanftnirpM5[M5Cba3M5Okaetirwf:oinY4Qba2Y4Nja>-)_(niamX4[j<[B9[E5.ba1|MOgacnirp(L5Mia(stup.OIT5Opa\\\\{)(niaM diov\\\\};)g4Hba5S7RoatnirP)--n;n;)sn3a<a(rof\\\\{)n tni,s tsnoc gnirtS(f diov\\\\{noitacilppA:RQ ssalc[\\\\{4&ha@(tnirp#6diaohtem06x23k+?a*3axam diov;oidts.dts tropmiz4\\\\{kaenil-etirw39lva(,\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'s%\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'(gol.elosnoc;)\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'K3s[2cya\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\' nioj.)1+n(yarrA>-)n(=ff4kia!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\}54,1\\\\{.n3cja# qes-er(a9dba&l5rba!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'9k$3lo3r33tla1% ecalper.S4l(3coWgsarts(# pam(]YALPSIDq6cua!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\".NOISIVID ERUDECORPU3kma.RQ .DI-MARG~3oE3dnaNOITACIFITNED\\\\{=dsa[tac-yzal(s[qesod(n6apa!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\");\\\\}\\\\}!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\");\\\\}/****/e3a\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"),s[99999],*q=s;int main()\\\\{int n,m;for(;*p;)\\\\{n=(*p-5)%92+(p[1]-5)%92*87;p+=2;if(n>3999)for(m=(*p++-5)%92+6;m--;q++)*q=q[4000-n];else for(;n--;)*q++=*p++;\\\\}puts(s);return 0;\\\\}\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\");gsub(/!/,\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\",s);for(print\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"define void f(n)\\\\{\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"00g,\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";for(m=1;m<256;m*=2)\\\\{\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"00g,4,:\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";if(n/m%2)\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"4+\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\",\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";\\\\};\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"4,:,\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\}\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"389**6+44*6+00p45*,\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";++j<=length(s);print\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"f(\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"n\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\");\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\")for(n=9;substr(s,j,1)!=sprintf(\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"%c\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\",++n););s=\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"4,:,\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";split(\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"145 160 17 17 17 23 252 141 0 46 125 231 229 231 250 151 243 243 243 231 231 207 159 63 4 231 249 255 191 22\"\"),\"& VbLf &\"(\"\"5 17 127 206 103 51 57 152 37 255 57 204 230 103 48 79 159 159 151 252 231 51 51 57 193 47 249 204 230 102 115 4 251 190 249 243 207 57 206 115 158 9 231 57 156 206 102 9 193 48 96 22 236\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\",a);for(i in a)\\\\{s=s 0;for(c=a[i]+0;c;c--)s=s\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"1+\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\"\"\\\\\\\\\\\"\";s=s\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\",\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";\\\\}print s\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"@\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\nquit\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\}\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\")');\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";FORiTO UPBtDO INTn:=ABSt[i];print(REPR(50+n%64)+c+R"));
$write("%s",("EPR(50+n%8MOD8)+c+REPR(50+nMOD8)+b+\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"J\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"+a)OD\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\"\");end;\\\"\")\\nsys.exit 0}\"\")]]></xsl:template></xsl:stylesheet>\":s=\"   \":For i=0To 7:s &=Chr(32-(Asc(c)>>7-i And 1)*23):Next:System.Console.Write(s &n &Chr(9)&n &\"  \"):Next:System.Console.Write(n &n &n):End Sub:End Module"));
end endmodule