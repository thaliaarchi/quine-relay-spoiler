module QR;initial begin $write("%s",("let s=(\"Module QR:Sub Main():Dim s,n,i,c As Object:n=Chr(10):For Each c in\\\"<?xml version='1.0'?><?xml-stylesheet type='text/xsl'href='QR.xslt'?><xsl:stylesheet version='1.0' xmlns:xsl='http://www.w3.org/1999/XSL/Transform'><xsl:output method='text'/><xsl:template match='/'><![CDATA[sub f(s$,n)print(s$);:for i=1to n print(\\\"\\\"\\\\\\\\\\\"\\\");:next:end sub:f(\\\"\\\"write,format=\\\\\\\"\\\"%s%s%s%s%s\\\\\\\"\\\",\\\\n(\\\\\\\"\\\"\\\"\\\",2):f(\\\"\\\"write{-}{txt}{echo -E $'(\\\"\\\",1):f(\\\"\\\"\\\\\\\"\\\"with Ada.Text_Io;procedure qr is begin Ada.Text_Io.Put(\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"interp:library\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"afnix-sio\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans O(n)\\\"\\\",2):f(\\\"\\\"{trans o(afnix:sio:OutputTe"));
$write("%s",("rm)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"o:write(Byte(+ 128 n))\\\"\\\",2):f(\\\"\\\"}\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans f(v n)\\\"\\\",2):f(\\\"\\\"{\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"O(+(/ n 64)107)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"O(n:mod 64)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"O v\\\"\\\",2):f(\\\"\\\"}\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans D(n)\\\"\\\",2):f(\\\"\\\"{if(< n 4)\\\"\\\",2):f(\\\"\\\"{f(+(* 6 n)9)48\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{if(n:odd-p)\\\"\\\",2):f(\\\"\\\"{D(- n 3)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 27 48\\\"\\\",9):f"));
$write("%s",("(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 36 11\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{D(/ n 2)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 21 48\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 48 20\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans S\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"STRINGz:=REPR226+REPR153,a:=z+REPR166,b:=a+\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"2\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"+z+REPR160,c:=b+\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"8\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"+z+REPR165,t:=\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"#include<iostream>\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\""));
$write("%s",("\\\"\\\\\\\"\\\"+REPR(10)+\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"int\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"+REPR(32)+\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"main()\\\"\\\",2):f(\\\"\\\"{puts(\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"class QR\\\"\\\",2):f(\\\"\\\"{public static void main(String[]a)\\\"\\\",2):f(\\\"\\\"{a=(\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"write(\\\"\\\",4):f(\\\"\\\"'implement main0()=print(^1^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"BEGIN\\\"\\\",2):f(\\\"\\\"{print(^3^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"echo ^1^\\\"\\\",4):f(\\\"\\\"'f(s)\\\"\\\",2):f(\\\"\\\"{System.out.print(s);\\\"\\\",2):f(\\\"\\\"}s=^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\"));
$write("%s",("\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"389**6+44*6+00p45*,^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";for(c:(^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"#include<stdio.h>^8^nchar*p=(^15^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"Ra#include<iostream>^16^nint main()\\\"\\\",2):f(\\\"\\\"{std::cout<<(^31^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"class Program\\\"\\\",2):f(\\\"\\\"{public static void M83abbSystem.Console.Write(^63^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"Quine Relay Coffee.^64^n^64^nIngredients.^64^n^63^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9"));
$write("%s",("):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");for(int i=9;i++<126;)[3pva$^63^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",2):f(\\\"\\\"{i\\\"\\\",2):f(\\\"\\\"} g caffeine \\\"\\\",2):f(\\\"\\\"{i\\\"\\\",2):f(\\\"\\\"}I3b54rja^64^nMethodv4f#aeach(char c in(^63^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")))^127^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")^127^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^32^[2al3dp3c[2cs3c,3l[2k@3kqa^31^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")s rts(ecalper.h3eja^127^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f"));
$write("%s",("(\\\"\\\"\\\\\\\"\\\"     53c4a SUTATS(egassem^127^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"rts(nltnirp(])]^127^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\".NUR POTSu4cba.C3dh3dX3bba[65bX4df5lp3lna\\\"\\\",2):f(\\\"\\\"})1(f\\\"\\\",2):f(\\\"\\\"{#\\\"\\\",2):f(\\\"\\\"};)06xt3dba;+3noa3(f\\\"\\\",2):f(\\\"\\\"{#qp]\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"};)0,#3rv3rR3sv3mba723284-fa(f;)1q5.ba.>4[ga#(f;)3P6[=43ba7=4.<4[<4[<4[v3gJ=d=4[73++>u?4[73xda,43?4[?43ma^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"' D ; EYB RCo8[.6[?4;ba5qB/daDNE&6[&6[&6[8Emca AL9"));
$write("%s",("[)6[)6[v3oeaPOTS^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'6[^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'6[^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'6[M9pL9[(6[(6[v3moaRQ margorp dne16[16[16[v3lbaST9[&6[&6[JQ[~6[?4Nb"));
$write("%s",("a4~6[~6[~6[~6>ba&g=[$6[$6[.@neaPOOL|N[,6[4@[>Xp>4[#6[#6[#6[#6[#6[#6\\\"\\\",2):f(\\\"\\\"}da&,)l=[^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'6[^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'6[eUnga. TNUO9@[,6[,6[83nearahc1G[)6[)6[R9ogaB OD 0hU[-6[-6[%No33)$6[$6[%NBca)Av=[&6[&6[HQoCQ[^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\""));
$write("%s",("\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'6[p=[v3npaEUNITNOC      0z41ba0y4.ba1>7[>7[>7[~Enf;[&6[&6[wEoRA[^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'6[^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'6[RAsba.)6[)6[)6[@4mja1=I 01 OD-6[-6[-6[C@neaA PU*6[*6[*6[v3:~6[~6[:OBxa;TIUQ;)s(maertSesolC;))T4[96[?4:ca11Y9/fatiuqnq41ca82p;[57[57[?4jda932A4.172"));
$write("%s",("ca65m4/i<[27[gC<ba9D?/maetalpmetdne.>72da215>7[>7[>7[?4kca007?/ca\\\"\\\",2):f(\\\"\\\"};^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'6[^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'6[?4;ca21A4/l41ba0j4[ha#(f;)34SA0batX6[=8[yE;ca64>HX>8[cCkda283m4[x5[v9gca5857/%a315133A71/129@31916G21661421553/:9[\\\"\\\",2):f(\\\"\\\"{;[?4:da429\\\"\\\",2):f(\\\"\\\"{;[b9[\\\"\\\",2):f(\\\"\\\"{;[x5[4Ewba0Q?0ra%%%%\\\"\\\",2):f(\\\"\\\"}*+1%%%%811 -%R2ca04"));
$write("%s",(";D/;6[T8[x5[j4Fca16/=0haj:+1 j@w?[W@[cW;ba4AD0D8[b;[x5[b;Gba8W@0baww9[W:[?4:ca13;T0>8[W:[x5[x5Gca99l4WU:[U:[?4mda818U:[<8[U:[x5[57wca05l4.baWv9[V:[KX;ca03=8[=8[V:[x5[KXw/?/ba\\\"\\\",2):f(\\\"\\\"{u9[U:[?4:da097<8[<8[3Xis=0bann41da364\\\"\\\",2):f(\\\"\\\"{5[*6[%>[x5[x5[x5[j4(ba9[>/X>[=@[8H;ba3=@[;8[T:[x5[x5[x5[x5[x5[j49da431l4.wa)(esolc.z;)][etyb sa)^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'f>[F?[?4:ba586/#6[#6[#6[#6mfa2200uq41da806-=[-=[F?[x5[x5[x5[x5[x5[x5[x5[x5[x5[x5[m4[x5[x5[x5[x5[x5[x5[x5[x5[x5[x5[x5[x5[m4[x5[x5[x5[x5[x5[x5[x5[x5[x5[x5[x5[x5[m4[x5[x5[x5[x5[x5[j4#ea2181m4.ba^1^\\\"\\\",4):"));
$write("%s",("f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'23(ba7@45ba7=4.da,43?4[fa(f;)5#6[#6[#6[#6Aba,%6[%6[%6[E9[#6[#6[#6~ba!m41ba6m4/ca~~37[37[37[S:[#6[#6[#6~ea(rt.(6[(6[(6[H9[#6[#6[#6~ba)BA[v3cda\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"};p4[SBfdadnes4[s4gra~~~~PUEVIGESAELPnr3ala~~1,TUODAERw3a:4[:4i$a(etirw;\\\"\\\",2):f(\\\"\\\"};u=:c;))652%%%%)u-c((||54[54ida#-<u4[u4ida||i15[15lhaBUS1,ODz4[^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'8pka"));
$write("%s",(")3/4%%%%i(g:c4;[04jr;[r;wPa2=:/t;2%%%%t+2*u=:u\\\"\\\",2):f(\\\"\\\"{od7 ot0 yreve;i-=:u;1=:+i\\\"\\\",2):f(\\\"\\\"{od))1(evom(dro=:t elihw?s;)s*z9[L;ny9[y9uz4[z4i0Adladohtem dne.s3dganrutern3dCaV);gnirtS/gnal/avajL(nltnirp/maertStnirP/oi/avaj lautrivekovniJ3d25[25i[2cib\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"};0=q;)]q[c=z(tnirp.tuo.metsyS;)0(tArahc.y+z=]++n[c;y:]q[c?n<q=y\\\"\\\",2):f(\\\"\\\"{)0>2%%%%++i(fi;48%%%%)31-)i>3c&as(+87*q=q\\\"\\\",2):f(\\\"\\\"{);22212<i;(rof;n)rahc(+O5[O5q[2k.4[.4%oa=]n[c);621<n++z6aqa0=q,0=n,0=i tni;R4[R4%oc6ahi4asdRbQeelxfvfXk8f<bedRbzk/2;agb-a|dzdxd8fGb8aqeRdYd5a\\\"\\\",2):f(\\\"\\\"{b2b4i;agb-epb>aqeRdHa>aJaRaAdteFbae:b6aOa5aaczg\\\"\\\",2):f(\\\"\\\"{fyb9a2*4aLa7a;a4a<a=hamkdxd;aNa?c6a|eebHaFaIaebzeJaeb9a/a6a2dQbUe-f2a-f9a2*5d6cRbC3gSc-f/aof0f8fQ"));
$write("%s",("g5a*h5e/,2e6aRa;d/NMfx*5h;aTapc4aLcEehiof6amc9lsbHg=,=fybxcxc>aGaUeAa2a6aZf7a6a@a1a:a?aMbKaKa6a?e:aA,2a?a@fMbAfGa>a:bXfYl;f\\\"\\\",2):f(\\\"\\\"{bHa4atc2iNa+bqj3bl\\\"\\\",2):f(\\\"\\\"}EcH=JaMa\\\"\\\",2):f(\\\"\\\"}bJa41Ec-bJaJaUa-bJaMdJa8bTaNa;a8b;;Ka\\\"\\\",2):f(\\\"\\\"}MepTaqjXyOaSa+z+b9bKa\\\"\\\",2):f(\\\"\\\"}M6*Ta\\\"\\\",2):f(\\\"\\\"}M\\\"\\\",2):f(\\\"\\\"}MepNa+b\\\"\\\",2):f(\\\"\\\"}qJaLaJa8bh7Nal4c#a8bNa+b4bNa+b:b+b<Uqj<Uqj\\\"\\\",2):f(\\\"\\\"}bJaHa#3cca\\\"\\\",2):f(\\\"\\\"}qm3a+aFdTF;a8bLt:aUa:aTaNadi9f7fAl4a*psbsb2be3^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'madiDa-a|b7E-aH6asaMSUe>auj1aKaKa?a@f*6cia1asbobdg06csasbHg*b-a/bxcHa|f"));
$write("%s",("e+e3c$b\\\"\\\",2):f(\\\"\\\"}b1aVg1aTfXf\\\"\\\",2):f(\\\"\\\"{bHae+8f-e:a:a\\\"\\\",2):f(\\\"\\\"}bHaYfJa\\\"\\\",2):f(\\\"\\\"}b5aAdte@aXfqie+xcpb7anb2b:b1a2f-j@d<f6aNjxcHa>aIfGfVj-a;fqi-fHamcdg9\\\\\\\"\\\"),\\\\n(\\\\\\\"\\\"f|fe+ze6g-fHaLj2=1ba01=.eb;a/aah<b=avh<apb/a2hnbyC7b:b1a/aah/adgbgFami|b1aGa3b:b1azhHae+HaUeniCe|bxc3b0a:b1aIa|bzeJa|j6biaQb-f@gmcn4awa-a5m*c3bxdUe=a-a?aev9ai3eraJg7apbwyVgTgRgPg9m3hCaAd9NPcgfvfxbydzb7awy*k|kMa5m*cEc,dJa>a2a:b6afjykMa?aev\\\"\\\",2):f(\\\"\\\"}i+cJh6a13eu3a[aH,+bvbng/a2h=aXhRalbOaCdlbOa4q=YNaXh1kDh7b5aLj8fwbijUe2bAdtl6F-bhcZmRjRjPo0c/bxd+h\\\"\\\",2):f(\\\"\\\"}hUi:@aea6a2bb@gocGW6avn2a5a3af@Zf3hRk6twjDhBhVmHa1dmd9h8f1k<kHa:e1k<k+l<b3bxd6a*h6k=hzl:uShxbziacPa;a,b<hQtfbpbE.kvZb<wnbNfajYiEc,d?azjIkahGktj<b<b<b3j:b\\\"\\\",2):f(\\\"\\\"}j<b<b,c8j5j<M8jEa0n3bDduk:i9a7blg-a5b|:,c8j=a9a7"));
$write("%s",("bcuq3e13eca0j13ceaIuxkA3c/3ggaJb7bCf#3coauj@a@aEj9ag*xb)3amaShjkVi5k,c8ji3a/a-a+bNg.bLg,c8jsb8fJjQk;k9i1jCa9i6aJjQkQjtj@6akaHjPksk<bzeVDceaHaZfM5cca,k53c/a;k9k3a6a<bShIiS=2b2a2a69Nj3kqiwbij8fTgnc:eUAa=aubzh5a=f=anbNjybnk5a,bJa6a7b5a8gwbijHa:e-b9a9b9aYjNjWf>am3awa@a@aNjWfTg:a|b9a0b9aTgUCaAa>e|b3g9bJa0bNjWf-b9aYj9aCaAaJa9bNjnbJa6a|b5a,b8f:e-b5aQmtb-aY;a$aPokPdi69Wf8bAd5h-a69*b5s-a69Wf7s3hlbPokPXb;d/g/bxd6a-b9a8b9a7bJcJayb>a/=Sh>aJa*c@dxc?b,bto>aJa-b8lteUeTg5R5aDc.G:atcJaub5aEc.G?a6F-b9gI7akaQjEk3amd9h^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'7g7cOkMkpb;awbijplVmWSsF49jN@0kPFcW"));
$write("%s",("lrlDmjn3lsnynpnj./n3z;03z2G\\\"\\\",2):f(\\\"\\\"{pXn*b@w*,+=nx-KC/h-C/bx*3U3t7\\\"\\\",2):f(\\\"\\\"{*G,f,ar+Ribip@Lf,5bZa>aEaUgf,,=n-vl1bQw6t@z*hwC7bCaKnBao3hbYK;0Wy5pTan@CoAaYaI|bA;uDaeq6bCa;0|bxpcpEo3xBpCiDaoE,bgb66,bfbkbLUd8-pQ*Eafi\\\"\\\",2):f(\\\"\\\"}5c7gPzfru3|GP7r9>ak\\\"\\\",2):f(\\\"\\\"}hbSaYaRpEa1bhbOwgVn*uopzUsS\\\"\\\",2):f(\\\"\\\"{ZpILYa>PT*h,i9q<AyM<avmIaqybXaDyttgMb/yob/I,Eo@ayb\\\"\\\",2):f(\\\"\\\"{bhcu21pazib,dgbhg4Thgsz/b=aV>yb6wxdp6b2:sGs9b8w<4FatbCaybHA\\\"\\\",2):f(\\\"\\\"}brY7Vr?C,I4,bdrXnIu4<Qan=Daib+bB>Cs,wl:TYQ=ecax?=TadvjxeTE5dsDaSnkpJz1K9CZp7AUad,-pG0@L.BlrDnssdCeq-08pU0Vs+t0<PnHMyb\\\"\\\",2):f(\\\"\\\"{b?sG22bqHOAFtQnPA*bhikN:Yib3oZo9Czb\\\"\\\",2):f(\\\"\\\"}O\\\"\\\",2):f(\\\"\\\"}bFrY-L*i9VahbNaam7Ugr2b4tabHun-RWt1e*W7n/ypibBah/\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"{@yfHFt7bzzP>nv@a22az.sgkR*BaNaTF4Imjy"));
$write("%s",("J/@j:T*c7Aagw?awbxbqHfbvs-b?nsqehY3?nnx;nLnZX//;:YaCo\\\"\\\",2):f(\\\"\\\"}-f||XCo=.t-4QZwG8Dy>av3hbxqwQ1buQf,+*@qqQf,y1OaBt,7ShroJ2YheT9\\\"\\\",2):f(\\\"\\\"}:S@tFJlbYPLI5xAO>am/Wa;6jb*bUsy\\\"\\\",2):f(\\\"\\\"{>a/KOacNu?0bu>wb8\\\"\\\",2):f(\\\"\\\"{@?Qsg.%3c>d>*<PYNVmWSf@;YxHfN@O-\\\"\\\",2):f(\\\"\\\"}>aShro\\\"\\\",2):f(\\\"\\\"{uCQeTDa/10bZSZAroIGSaDaz29\\\"\\\",2):f(\\\"\\\"}e8;|QaFatbCSybRTMnz2f,,vf,AO;zM/g-jb3mgbcxCaNaM/g-VOUa7M?n6qSa:uFOnsEais,bC/OVTn2b0v,bOVTnj,>PzbQnmbgOU\\\"\\\",2):f(\\\"\\\"}g-ZV/K6b,bZaBF=ankiqXaMt>aIJ/O-\\\"\\\",2):f(\\\"\\\"},GU\\\"\\\",2):f(\\\"\\\"}aoS|MnH?f,djUs4bSaQ30wvT6bOaf,jOMnvb6b6|v,f,;qPPSnJ;BF>aPaF5Ua-zQt9*|:@-i2Pajb@a3ofb9b?Wj|NaQ+M/vs.bSaM*jbDavsy\\\"\\\",2):f(\\\"\\\"{M*<30bgb?NW9a^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\","));
$write("%s",("4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'cfb9b3b0bgbxq|2=a6N4Ngbjbm\\\"\\\",2):f(\\\"\\\"}Pa-bvb=:jbMMjz2bnQd-y|*pzN.U7b0o935bjSP\\\"\\\",2):f(\\\"\\\"{1IKnJx:7vshbNaCaRROZMP0b8=6=?W=aM7Aa+,hbP2DaCn4ThbA<MPOkP\\\"\\\",2):f(\\\"\\\"}q6CLpm4blb3bjohb,kqzg-y>=aKHzb-pMPOky>YKb\\\"\\\",2):f(\\\"\\\"}9Mhb,kDa5Mv1FYFtn0QaDaj+JwhbF5OahbRaUwhbOkl4cXaqp4b5bVJDa+4xbLSK*gbdw2bDaMUZaApDpab89mpctBaibmbGhdQsPDa,oyYlt5M|<ZlDogp35lb9OBio=j-=b4bAtzb1,=a?UqpL5l:;wi-<TZa6TcqbbeJ>-<a=aLvKBU-5@BU70hbhb0b\\\"\\\",2):f(\\\"\\\"{6SE+<:=e=ZC\\\"\\\",2):f(\\\"\\\"}5=a5Ba-\\\"\\\",2):f(\\\"\\\"{*IpQn+b:Z3=ySZa8\\\"\\\",2):f(\\\"\\\"}5,DtBq=aJxNkTaGa=O<aTa4wYaHyhbVaB>d+84tb$4a,a,bn5;<Q+2b2-t4\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}o,3oYaXa6848Fa>sBa5bW6i)3drbibItpzFv3-Vqul61GSTa\\\"\\\",2"));
$write("%s",("):f(\\\"\\\"{2v;a,\\\"\\\",2):f(\\\"\\\"}yGOetNR3bjom+rqvvXy+*9t3r@v+djoib@L3oBaNa8\\\"\\\",2):f(\\\"\\\"{m+,bI@,vebm+Qq+**b|d5-HAvbQq1pVTIW~DcQcnd43avzt2661DaR/O|ERm.s4I>Xnp8gbNxM*Uav5H9P0Oam=0*8-cU2bu2RtPDkbUxb0-<>rLVLRC=6wgb\\\"\\\",2):f(\\\"\\\"{9\\\"\\\",2):f(\\\"\\\"{b8tZal0Lg0bZS8S2|mIOvebWT=:OA,DMt8r@.>|AO0*+bRq/N|+GadxrqU|2b:uX6./QD>aybOK<aSht-BA>adVbzU8,btTZ+d8@4?WNAHShAG@,DNkKCPRtuBR3/Rv:7xbdbGtgbOyub0bn=CQzLbwWY\\\"\\\",2):f(\\\"\\\"}bUp2*Ga=Okqf4aya|GetEaXsU.Q1,kSh.9n-OT,sC9azdWaKH-p6hbA7bK*hxgmf+*<T?I=X.1bp0A,1Q-Lu/\\\"\\\",2):f(\\\"\\\"}ydVVFj|VyNaP=mb9bsvzOVObzhbN4ZaUu,b1bXaM;-Fo?\\\"\\\",2):f(\\\"\\\"}bg,Q*zpgxSaZGEq<afba+9b|d3r@v*/rq-FdJ+F\\\"\\\",2):f(\\\"\\\"}FCv6s*:M|ub0bsv*:S.6EfbVM2GZVbbIwPwwb|,3uY-bbNaRarycx<a3o\\\"\\\",2):f(\\\"\\\"{q\\\"\\\",2):f(\\\"\\\"{Kdwnu*bCQR20z9UubAHab+yLrhbPfuVIrD\\\"\\\",2):f(\\\"\\\"}C|84s|@a"));
$write("%s",("a5;U02DrZr7\\\"\\\",2):f(\\\"\\\"}TsVJSh.9;2Z/9tRyS\\\"\\\",2):f(\\\"\\\"}Er/Bk>;|xbG23o@+=aKONA44+JcKe+aR=1bvb;zN?,b32Va0*0z;|vv0*PVqHtyoC0b\\\"\\\",2):f(\\\"\\\"{bjDeuawbZs;9SadJX6x*O0|CJK\\\"\\\",2):f(\\\"\\\"}3eVbdwCaub0behs|P2x,+b;2is@yk>,bd;nLFYEaw>T\\\"\\\",2):f(\\\"\\\"}D504>P,Bk\\\"\\\",2):f(\\\"\\\"{pZAa6xT9N+j/H*fC/b-KJSv=UsQ|-/qH?pmR.b06>\\\"\\\",2):f(\\\"\\\"}Na|>gbG23bSye2qH\\\"\\\",2):f(\\\"\\\"}T1uGSSaTnvxM@\\\"\\\",2):f(\\\"\\\"}8Sa=\\\"\\\",2):f(\\\"\\\"}o+7b\\\"\\\",2):f(\\\"\\\"}8m4u3e0*bybEah-,bRaTaNH2r5bpTm3cutb\\\"\\\",2):f(\\\"\\\"{3akaKB?a>P|,Vwo3aca|*/3itbI1kb/N61Pn\\\"\\\",2):f(\\\"\\\"}8Qybs3o1b0lkN:YD,I1Zp\\\"\\\",2):f(\\\"\\\"}ur9+Exq77In7twQZa?4Oa\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{Yu1HgbYa-zA5gk.dybE5vo-pHy7|jb*,xM6wSnJ2P*;ge^127^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^32^[2fha\\\"\\\",2):f(\\\"\\\"})3(f"));
$write("%s",("\\\"\\\",2):f(\\\"\\\"{#v3rga(f;)0,73-)cG,/TaS;?acb3-1b3o?=i,WaWazO?=RDyo>o.bHXL+9Z9x.b@.kb<a7b\\\"\\\",2):f(\\\"\\\"{v,5ub*=JrxZ-bnL<v/bXt5b9NRNUaZrsv6x3NK\\\"\\\",2):f(\\\"\\\"}<-s;5PZ/TndbcYIqmj*bdVmV5b+qxtCIab<-uEur/bNZ7VxEUs7+dqNw\\\"\\\",2):f(\\\"\\\"}Nh7/BJDFa0+jpS|:|Eag,=WK6=alFKB?a02.6v@2b:1eu8\\\"\\\",2):f(\\\"\\\"{pso=Ua|15b4oEb|d6v7K/@.WNa+2/behf2ML-:0bitNaAaHSNLRtGsEl-r\\\"\\\",2):f(\\\"\\\"{63be,dpBatqu1s1Q\\\"\\\",2):f(\\\"\\\"}wBgMZ6Way2P=TaCE>qj:otZt7TBajb\\\"\\\",2):f(\\\"\\\"{bUs3BZq*s0bC|84Fa*3,bD<<zPa@a7bhs2bb*8?<a@y+d*=JKUsY0a,Y7;z/bER/x2bOaJzibSaFxy?*mBxspmbUaEasy33i4cQ|;Wa7;DNgJHyQx:=vRgbn<2DtbN3-:ibibm|ArVEaj=/-dCxg*c1Rptvibibo|lrBAUJNY2b1GU*p\\\"\\\",2):f(\\\"\\\"{y+3rEx8Y6wXaqx0vPV+6$6aAavbFaUa;Tuv1bLgbptzDvtTNEtztqeu8\\\"\\\",2):f(\\\"\\\"{YnGa:R+bUpr*6hQa?5=5Vagv4.7;sIaRbuq1bjxG*G0pZAafSztgvuBVT-i\\\"\\\",2):"));
$write("%s",("f(\\\"\\\"}-c9Wqbb9bamSarqZXGoG\\\"\\\",2):f(\\\"\\\"{CaQX6b,bzNK\\\"\\\",2):f(\\\"\\\"}QabbK7FyOY:4<wGaq-czW82b4<mx2VWpK77x4<|Lh/dD;R4/\\\"\\\",2):f(\\\"\\\"}-Wp+qSa|8Ga:R,U./8p@nP70wt106i\\\"\\\",2):f(\\\"\\\"}QahbaFyC7bP\\\"\\\",2):f(\\\"\\\"}vo<a3oM2>aPae3a=aQ-xbtb3BS\\\"\\\",2):f(\\\"\\\"}/1;1MUlq7xtq-b2EC\\\"\\\",2):f(\\\"\\\"{bwWYGzA\\\"\\\",2):f(\\\"\\\"}NakrRvRx7EF|7bl>x9+q(6amcQaAvr8AvhsX:,UU>LlF*Aqptgve1B>55bv/bNaDNRa=ambI@Ya99?o5xouw6*s0bt6EalbV/MIfbkbTuGa<WP.dodSVa?oYa\\\"\\\",2):f(\\\"\\\"{uLUAacQXaV/OaDN\\\"\\\",2):f(\\\"\\\"}b*40b7tw6HOYa/>*rGa<Wx7SabN,ba089ttjCGa<W89BrdI.Bvb99Ws6Cip=/jd.EldZ6*b,?;3aub;;Way2=ajpbbCIQFjxhbLS/@.Vcqq?i4eb\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}dJLr8\\\"\\\",2):f(\\\"\\\"}lbF*UamI::q9l>2bQ|*=MtjSmIg-+*?aPAwb;*zzzo>C184blbmyl,54Q\\\"\\\",2):f(\\\"\\\"}5*kCCs7\\\"\\\",2):f(\\\"\\\"{=boc,bZa2qAD+*0*n.54qx+qAOlq/stq+\\\"\\\",2):f(\\\"\\"));
$write("%s",("\"{Qa4v2vcO2bmIrqPVe,qx+qrM7=P,WarPhM*q1boxyA5=;qfbdbxbySv=@S<vf-Q>PcnUZakoGadx1*:zj+dbUg5=?UfbaxgO4v\\\"\\\",2):f(\\\"\\\"}u2sy*Va20JS2bL*6zvsT,Vv;CVEpzw-+OY3AoJuDalqq7HXL+*O|bs*GQSR;3cia<-NawEI|M3e6b<a015qT\\\"\\\",2):f(\\\"\\\"{yAdb7h2bHvCNOqC:ecC:<vqHl\\\"\\\",2):f(\\\"\\\"},b1bBAI,2O+yX6,bFP1o5=uJkN:Y?aWqF*xbaKeJGaSYzpaJboh3fQg=eGCalq>CtvFF0vkbN43u6vQapm,Op6<Lr+DSAY1bhbx><Wi3a#ca,2bN4SaRTXaLS*:Na*b1*,?.b|X|i?a30-:mVJ3do/bxr<W\\\"\\\",2):f(\\\"\\\"{bQ.0Eeb2*-:;/EY2*-:=2FnBtZs1b*4R2AY1b:P|LN4Sar*TaHv<-L*QaMS<W\\\"\\\",2):f(\\\"\\\"{bBn/F\\\"\\\",2):f(\\\"\\\"{2pZAaDaDvrjWq3.|XOnE2CS<TMUgBiz2UH=W@zbtvRN|Xdj>amCzb0bb>?amOWDOK\\\"\\\",2):f(\\\"\\\"{bjbbb2OqHTu5Sat/B91or/9a/a-bt4Ou\\\"\\\",2):f(\\\"\\\"{bBas;-oqz2|C|9|3o:oUAnMup+gI4\\\"\\\",2):f(\\\"\\\"{b\\\"\\\",2):f(\\\"\\\"}wS-~6c[av>2UmyTHNa6|qj9<M?Bas;SayuCsO\\\"\\\",2):f(\\\"\\\"}hbTvM\\"));
$write("%s",("\"\\\",2):f(\\\"\\\"}|vVOtv*/vseb:26q0p9*ZqDS7b54@QmvkbkvivTa0,?G\\\"\\\",2):f(\\\"\\\"{bZa0C^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'H(ba7>Hv2Ivba72I.da,43?4[ha(f;)594A4.ia(ntnirpnt41da652t4.ba)T5[97[97[v3l@bAT@a3vQ1Rqdt2B>PZa/BY7w>\\\"\\\",2):f(\\\"\\\"{BFnNaKsvB=<B:;q0bEN?aUa5bF9uB=a:|,=|rz8Bp.Gjbx0h-m;-4bSN/m1Ex1y>amEbbYakgM+>yhb0b3Ldj-zR5@7Fti\\\"\\\",2):f(\\\"\\\"{PabbhcJxEfe-A9Yaj-=amb>y@zrWedfWeP<FxXaAzqjhcc6NT+;;;2IebShLryum1:\\\"\\\",2):f(\\\"\\\"}/155ibVa/5Fa5.|*jkubRa@L>aw5@v>/0bX+8Y5\\\"\\\",2):f(\\\"\\\"{Qabb.Y?a4bxQwb67+,On?7o\\\"\\\",2):f(\\\"\\\"}=/6CXa7U+q8/t1q7fbab\\\"\\\",2):f(\\\"\\\"}u-<WTao3/Rv:7xbSh87Z*Z@ybxb47m"));
$write("%s",("7Wa?6i.f?jtd:-thv*u,b,7OyJdXa<albDaU-|KSAEZE6:yRaUgr+EaybShQ=<Nfg5Ks0M,Y31u7U>a1Q9=<aVp,w?noIRqYaXa@P,DXTB*1*;jFOX*kbuq/bwDfoP.OX=apNlR=aDEXv;YxHiN49jNW2\\\"\\\",2):f(\\\"\\\"{bhMam*b=*1bmMHOn8iRCajk,b.bv4c,+ccbs|v>u:z2Q\\\"\\\",2):f(\\\"\\\"}.d@a|d8-V*h>bQ\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}jxvCTnXa3oybUU0vGyrvSqH/-bjbAag,+4Cpkghbn\\\"\\\",2):f(\\\"\\\"{7B04KIf,xbQaB:2bCvN/Qaz/s@a@jr1Na.bbYAa9bvCA1vvh/Y-oxmHMOyC3bFM3;qhRalbTPwbpqZ:/;=aVaust7,;h/++N;A,j-Va9;84YPsK58tbGuvbnX?=tZ</fg?ARaTuv*2:n*sP2N@oLSCfSha;U@;=3be/$Y[v3bna1=aWU2txb+;Y:wFa~djkbIsyNa=;ib,uA4Yh</fg?|0;.;SaWaOaZag-j7\\\"\\\",2):f(\\\"\\\"{;TuPqHh\\\"\\\",2):f(\\\"\\\"}Cvbpq=;ib8riQEaxbuGW<f;Ra=;P0ErlqEasy:z9bi7,;h/=asye/-;db,8lbsvk0IYl7WaAa>|-r0@.@gJ|6zb:|Xn/gu7HGcrvWVadMwq65@y7\\\"\\\",2):f(\\\"\\\"{CQjb\\\"\\\",2):f(\\\"\\\"{9@Lxb1?rv@aNaW;u?M-dW3ofbq"));
$write("%s",("MgbaF-0QXD3Pav*/b@aPf>t.bC=@r6bRH.bNa+ba>-tY-0bAy:z+>s|NaBwQ=jt7zVsNOBULE9ktI2b1R4bzbGFc|5q1bEaA4@Sc\\\"\\\",2):f(\\\"\\\"{d<gDo5Mcr/g,d:=1:QGU?65Vi;rQ0:/ZauO\\\"\\\",2):f(\\\"\\\"{**bS3s105pmv3hb.bC,\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}jxyyCa3./-=Y+uGu,bzJ*QVa;IERn22|qH:;9bwbur/b=a<a2LI9Wa-o-/SaAam7g2ufj6VENa+*WaWausZ6:ne7TPc7mh3iDa=af9gyr?Dy;2c*1BhkZavbhbvT6b;qDar,E5FEazFE,rL5e/TP0*ushcDassLE/gqxRa?arP0pYau2?3|;5V+CAK/8UasCRa1bIdDaa,Efjb/NfUXJ-r\\\"\\\",2):f(\\\"\\\"{60+Dwd-Na9-T/0blfMb@aPa7=>atOmvb6zbv*+b\\\"\\\",2):f(\\\"\\\"}bTaJunv*,9kk\\\"\\\",2):f(\\\"\\\"{8WT,YPn0PS.babPaVo|,jRu,efwa5f-cUawv6bi7mR@akpiFv=Usg9>-.sY/|LO|<\\\"\\\",2):f(\\\"\\\"{jbubDp1Yxbd\\\"\\\",2):f(\\\"\\\"}Q@O@>@@aOyJdO|VGhMQ*gx,udwlrTpbz=88bV*m1Ga=OxbcB/\\\"\\\",2):f(\\\"\\\"{bqdb2ODv<NmpN\\\"\\\",2):f(\\\"\\\"}L\\\"\\\",2):f(\\\"\\\"}LwPPqAg?wbe,y1r9JUSh=U\\\"\\\","));
$write("%s",("2):f(\\\"\\\"{b,bzqcoM|5btvkb3vo:<-db2OTZldUadbO.mo:\\\"\\\",2):f(\\\"\\\"{kbNO?oC\\\"\\\",2):f(\\\"\\\"{Aobb<a\\\"\\\",2):f(\\\"\\\"}b?a4B2B6V4V|+lp4yS|=a@+aj|6and8b.B,B>Vco5+3rit@WibE6zL@wUxkoAC/gS|2:\\\"\\\",2):f(\\\"\\\"{7iq>PDNYaY7Q2\\\"\\\",2):f(\\\"\\\"{YG5E5HvGz*dcB1VS3Y3;UKI?7-tvtXajbc?x*h-nrEaBae+sTnBd-lMB*Na1vnrcoXF3btv4b</QA:Pyb6bYjBa,b\\\"\\\",2):f(\\\"\\\"}32x*4Oaz>1bXajbX77KEEM|\\\"\\\",2):f(\\\"\\\"}3oANnHA+blB-rybsTgVzS=:b7v3at.bjr\\\"\\\",2):f(\\\"\\\"}bR*7Ku84J,9@ont,D6FibTKj6MwLxsDxbab>s4exEjCRyMvbbAaX:Wn=aY/pNQsMUSa44q71>r6a1a\\\"\\\",2):f(\\\"\\\"{bv*>qCgA.PUVa\\\"\\\",2):f(\\\"\\\"{1d9Gy,YSEg|+brqQQ\\\"\\\",2):f(\\\"\\\"}sCigr\\\"\\\",2):f(\\\"\\\"}bhbjt^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\""));
$write("%s",("\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'Ga/a;rUglDA|7sM\\\"\\\",2):f(\\\"\\\"{GPpEfUVqf,n;8-L2GyL2zbYw2CZEsC;3axdff3/;797h>..atCgbbbbv*c9?3QyXa6848F.LSi;lpAE>a\\\"\\\",2):f(\\\"\\\"}b02hbc>6-0CZajbCaotqr\\\"\\\",2):f(\\\"\\\"}t9bat7bhb7b+D>oab/KVymFWarEe*ZaupZCJ9|rZ=lDrhXaxb/NySehVFK|ERl,u3Aav,vGlDpmvbhbaoUakgu*HOj|sy.GhbtqSaeCPM@a\\\"\\\",2):f(\\\"\\\"{6+bBaebVmWSf@;YxHfN\\\"\\\",2):f(\\\"\\\"{Azbdubb1olbbb,v/-zbJd>aXVstZak\\\"\\\",2):f(\\\"\\\"}TuMtO.-\\\"\\\",2):f(\\\"\\\"}=a2|1<TnQad1.bT\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{b.;lb+b,pw5lbfCj.V/Aq1<AaLI?p1Q)3a&bj.9LVwE*j,e1qsKN+bz/oUBa\\\\\\\"\\\"),\\\\n(\\\\\\\"\\\"1GjAnuN.PqBzPq\\\"\\\",2):f(\\\"\\\"{bXHScBaQN+bBaZ\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{A.dHhO.r9Lp<alb\\\"\\\",2):f(\\\"\\\"}Ky|FFUa|sx1cbEa2|1<OajGv,jGjOZ6n\\\"\\\",2):f(\\\"\\\"}yz6\\\"\\\",2):f(\\\"\\\"{9bPaJD-t-*Zwc3iCaybV2C8*hC8*h=ak**b0b+bmCix"));
$write("%s",("bb7?NZ/8\\\"\\\",2):f(\\\"\\\"}UzpwQ5t/|@QkbMEhbnqg>CrboybG9a$dYa7;zb1bpNmo?atbDa3zsszblQ,x/=EaaxnMs;VaXaeT3v*,UatqxbHOD0OagwB=wb7o@w\\\"\\\",2):f(\\\"\\\"{6;1uEwsGa:4?9eh*umVi2PaPfwbj|@w\\\"\\\",2):f(\\\"\\\"{6H=3OI,4wecMs3;s/ibHSS1Uaehk8Sha;m1ysD1C|\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}NTjp\\\"\\\",2):f(\\\"\\\"{2\\\"\\\",2):f(\\\"\\\"{;qqn5/NR.XaArL27b=a9ZWp0vkqtbYaW8OYSYhbjvXQxZD05xRa.r41HO6s-rg94N//fCLE4Y<vxuv//BOz*5Q.Z\\\"\\\",2):f(\\\"\\\"{H4zqQahbfHr*Q*zpgxSaZGEq<aavQatot-zvLy9bGoTsZOD>ub2Re1aNr;P,oi2mwW@:ZD>ubtb4mMUFa;9UaapibxoZuSEgb4qm3e7t/1GS.s.I|L0bj.Va,U6zUp6oBZjR|bN+wNQaDv+bb**3=a.by4X5pz8K.VZaubT-UamV6x?Bmwap<s5qJ<C4<akbYaws0b,3d8y2Q\\\"\\\",2):f(\\\"\\\"}z;3o?aNO7;XskpXol0J;7uNYJI5bkbgy41syfbvo/BrPazAEbbT\\\"\\\",2):f(\\\"\\\"}hZ.BeD/tA1-h1oI/mbZaY0e:Y3Q*fPkbF:Z*Sh>wmjFXS+GauFr?.B0pm3RaSaIJSaeb91cu26Bz3bmjgbXa"));
$write("%s",("BceRFW?DSi+Edb|,5;6b?s=sbG\\\"\\\",2):f(\\\"\\\"{bYa0-kbNRZlE?wbzbYPfq8v?nbQrY0*tb6b|dkqCI?U?aRawqC/hMC/m4WaZbBa\\\"\\\",2):f(\\\"\\\"}s4NMI9bB1,ddb+C+bhUZaMM>aRp\\\"\\\",2):f(\\\"\\\"{K.sbbnimQh,JGN+CP4bQT19NO\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}jXW@NiKOZCnBr|Tp5;pLz833>MwDSa5bH.Aa1bq=sI\\\"\\\",2):f(\\\"\\\"{bcX-05-fbfbBUct5bCI8*:UcbVy@<cwj-DWfb>a0*n@XaQ58WVW3BdX8b90vV4NBa8b;<Xz2W+b-*Q0WaTMvxrL6<;PyuQps-fiXSyHRUg+,xr1+,<Ngt-bE6ShqySa=/R*JxN4*.Huw+.WCIHugbY|3bmxjba\\\"\\\",2):f(\\\"\\\"{ubjkbvLvcrFGJ;,bbzQ-cEybeNYa1\\\"\\\",2):f(\\\"\\\"}qpg*Crmj9bdb;6v3@.7slbtsefDrHS<-OycouBKj2GF\\\"\\\",2):f(\\\"\\\"{fbhVj|zbAamgzp7\\\"\\\",2):f(\\\"\\\"{KrzLLUlpssqsU\\\"\\\",2):f(\\\"\\\"}Oy<2;VwV.|7V+b=*fbzbK=J5|zFa>tUaLSNAdbzbeh/NlbQn8*Up+EjboAYjbw=r22\\\"\\\",2):f(\\\"\\\"}uzbZa74OnI|KutvO.bpvbNxf|WvT\\\"\\\",2):f(\\\"\\\"{u,ZatyV|cbDACa2CgwKBI|PuR42CXrjLVSc"));
$write("%s",("bQaKwL0hbCa/Kc;s;lMTp>qv>MvT-?acNwb2bE23b+b>afb8\\\"\\\",2):f(\\\"\\\"}3+tbqmC=HMKI2bOKS1CaDaDtabbrKOPauf2p+.j*A=bSz;k426l=@LZpzb+b=/wQCN3iDvhczJ99YaQwr?Ya5s3s:=i\\\"\\\",2):f(\\\"\\\"}hb4b3oRp>auEvb-bO|<a8bkb=NYPS6:Jp8y8C-Zb9kLSJn.bcbG8WwuDQaybd8.|6wabybU.abF:Taeh*Ts;>Sl,v*mswb5b-bB=5+8bZ7;0gbyb.bmblQiQPar,h/cbV0:sgtwbXJj60AlbN2Qq2Cipc?\\\"\\\",2):f(\\\"\\\"}liPV=cRub21LJZw=/6bEa?aGarSo>\\\"\\\",2):f(\\\"\\\"{b24wbdb9bGaYAib2GOxUqU3<j;PkbNBfQhBIw3;WnbbB4fSlb\\\"\\\",2):f(\\\"\\\"}5Y3-Ogb=,PHabn\\\"\\\",2):f(\\\"\\\"{bN1ubjlb,b02Rq8?24JGBwm:4t44g1/1\\\"\\\",2):f(\\\"\\\"{*V/azgbnv3.Zanq;qBaXs.b<4e4;w4NNEXzybS4Da.bM+B<pNc\\\"\\\",2):f(\\\"\\\"}dvxbrh\\\"\\\",2):f(\\\"\\\"}PavYuB1hbjbAp*:5babTHnxzts;uqShz@7R;2zO<a2b3\\\"\\\",2):f(\\\"\\\"}rCjxbbXa3wG,kOk2>P;?uBFNtb@2C3*soA3b:uW.7b4bGulsfr2Qkb+bXF9bYav3/bhihNg@hLe1x*VuUa|bUalbQwgAICO|@a"));
$write("%s",("bb+OE\\\"\\\",2):f(\\\"\\\"{CK>*P;,b\\\"\\\",2):f(\\\"\\\"{4*6vGfHv43BPa3o:-2bP;e\\\"\\\",2):f(\\\"\\\"}m3ktXaSG0bOa\\\"\\\",2):f(\\\"\\\"}k\\\"\\\",2):f(\\\"\\\"}-<jp-r*1uSadMVa26;<<\\\"\\\",2):f(\\\"\\\"}Q.DaMqCLc1I2P\\\"\\\",2):f(\\\"\\\"{kbEayu+*mP+*6|m1EjYnWnfb\\\"\\\",2):f(\\\"\\\"{b3t@albK.hvbAuo\\\"\\\",2):f(\\\"\\\"}y>aub@n<zaby*5xJrmqAa-/Q.61cbK5PHhbG8WHbv55K7Va/bP\\\"\\\",2):f(\\\"\\\"}M+kxg.Q9,bUs,b-*K,hb?a/ty>vt*sGt:|y*p1bb5y1I|bS|i;?GSLtb.bl0h5E5p6o,;s4b^127^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^32^[2fha\\\"\\\",2):f(\\\"\\\"})3(f\\\"\\\",2):f(\\\"\\\"{#v3rga(f;)0,73-c1-OmbwbeOcbPa0blbVmhPq5kLhDvH?a-bCaAsK5KNkbr3Lu<9Oa?aKO*sIOmdajxvVaPaa,kbbMHuwb3oebQA6q*szLDa/B5tvF|tl>.|61n<<x*O8KkpaocbOaQg\\\"\\\",2):f(\\\"\\\"}y\\\"\\\",2):f(\\\"\\\"}sM1EaQakbib<ah>*s3oe*fotb<zDaRaxdZFuvmO=aJ56b:2+:dbQg*rA9\\\"\\\",2):f(\\\"\\"));
$write("%s",("\"}uttaj0bfrfK6zI=6buvS.\\\"\\\",2):f(\\\"\\\"}bv*T|*blb=4Z\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}kNEfb=aF|\\\"\\\",2):f(\\\"\\\"}k..Hu<tQ7UacbKt\\\"\\\",2):f(\\\"\\\"{bw0qm:p4bmb\\\"\\\",2):f(\\\"\\\"}b>M/bm/|;Wyhb1bCaSazbPfxb<zs-@L*:NiFa1\\\"\\\",2):f(\\\"\\\"}=5gyR,Vy93z.j|nvDF1bt93bqH5bdqfiY2gNC;B0qFb@cbJnvb7bP<E*p+?xCr+bT*21VyWnyMBau,b/ubvy5M|b7oUa0b>a,bQmCLJKpLQGBt3bO6-bQm|yjo8/kbxMjbiv3DFtq=nuuwc\\\"\\\",2):f(\\\"\\\"}NitM@d,.SaQadb.o,xtbn*<8W|Pavb,bm1kFUCdbBa3bAnr?b/8bvb9bGy0*@ySEY\\\"\\\",2):f(\\\"\\\"{;1\\\"\\\",2):f(\\\"\\\"{1qvy|0*I1UCXa/9qs>yasXa=\\\"\\\",2):f(\\\"\\\"}y10b66|bv3|KGp6o6-vbS.WpDa\\\"\\\",2):f(\\\"\\\"{dbb9+U-W8cbVa2b/bsy*b1IAa*bbzh7|dh7-b;Bu,Zb1q/bQawbcqztZ\\\"\\\",2):f(\\\"\\\"{N4u:\\\"\\\",2):f(\\\"\\\"}bbD=;R4zbSak07@PoJ+sJU=qJv3m/?p\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"{dDi;-tb6jb-\\\"\\\",2):f(\\\"\\\"}Huj:6b,p@?jFkb3;yb30\\\"\\\",2):f(\\\"\\\"}:y1xD"));
$write("%s",("\\\"\\\",2):f(\\\"\\\"{b2.-w+ww7F=I3WaG3TaDfDokdgqiBZ*zzRaFa6b3b2K|bVy5b*hI|-b7bTal,1,TnmbTagbQC9two6ht:K7Wxlb*3XGyJZJqvWo+>?/Vna?L|OnZ\\\"\\\",2):f(\\\"\\\"{7;InGnEn8bG0*z/b\\\"\\\",2):f(\\\"\\\"}y?aubdbauzsC*AxR0dwCt+,6*I|lb?HppSaibuy>/</foXoLqebP\\\"\\\",2):f(\\\"\\\"{VEy1,?O?SEV5KHV\\\"\\\",2):f(\\\"\\\"{s8q8Ay8b\\\"\\\",2):f(\\\"\\\"{uE*\\\"\\\",2):f(\\\"\\\"{uP>ip-bAaCt<-9bkbybBazbwAhizHA;b3wHXvc\\\"\\\",2):f(\\\"\\\"}InSa\\\"\\\",2):f(\\\"\\\"{;F:D:b\\\"\\\",2):f(\\\"\\\"{d4mbh:tbSh|@z/hk|rH8Jwe*ffY3bbe-6w-d7=owTHlbNaQa1bGr6;J<gmitQmubr,EwnpAzQ0Ewm+9bq=Gt;8W;Wnfs=v9bBadb3bm@|bQpn*s|\\\"\\\",2):f(\\\"\\\"{9Qyf|-?8@6@aq=8H,wr\\\"\\\",2):f(\\\"\\\"{bCap1O>;H/b=/-bZCU?S?IxF:-0tqd10bb5@a0b\\\"\\\",2):f(\\\"\\\"{qZvcbR1,r@4/bn=<a5odbyb?ads/=cba?Grn\\\"\\\",2):f(\\\"\\\"}=aRa.sNgm+tb7bO?Ea2H-*nrjbjtH21>30Q3<a+b*B6bhbpo\\\"\\\",2):f(\\\"\\\"}b0\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"}"));
$write("%s",("\\\"\\\",2):f(\\\"\\\"}UwW<*dKnSEfiiDrFy\\\"\\\",2):f(\\\"\\\"}pFXaE62bFaZCQan,Ux8bWa@abo-/s7*,Ei2bGFEaAaQvasbbbr9bRambcb8xZa-F0bT45mDaOabpB@DaAaub*89b=agbCtV@jtAa4bpu\\\"\\\",2):f(\\\"\\\"}bZCk0/b\\\"\\\",2):f(\\\"\\\"}5Eqvlc9;BC*<aebxbCa19vbk2Qa4A3ou9Ba<aPsv*=/?aPa/bL*@agbabN4B>>CFa6<3=mb+t1?3/qv8bM45sFa=z8bWveb93jbU1Vat1r,cbRaarl3;n=z*Fh/+<tc7bzb+q7;CDvbfpo8fp7bd\\\"\\\",2):f(\\\"\\\"}D3Ca3b8DmCsq4buo2,5xwDxbIwiq8x+bs4a+0b,tg,qrubT11v2BShF74ad@h@@;gDQ1zbfbYa5b>abz-op,ty,:dsT1hBTa|b>CKCHDcb.bICXazp7bFa*mNaDaEa+3Fa6o2bD++bYaYa@aN4Vag>bz2CUCmd>a9byb*b*bFajEO?*bkbnE<-SvNa6hc9.bYySan->aKjSacb=abC5bh=Z*lbHd,rRa7b\\\"\\\",2):f(\\\"\\\"}bAa?DiqmbyC;1abCBzcVa7>2CaqCa+bCa\\\"\\\",2):f(\\\"\\\"{v*-Ryco>sWaKr@aKjd;|;0wtb?CY-U-f;1>?elbz,Pa?aCaibdqbqDv@ajk*mOafbU-;CRaybgbbDCnhb0ozb;rb|=aj:?oPv1,|*7bx0,bi+Xo|b1<6r;rcdVaFa"));
$write("%s",("U@\\\"\\\",2):f(\\\"\\\"}lW=c@WA0vSafb<acb/zYav>i9,4?\\\"\\\",2):f(\\\"\\\"}<a*b-\\\"\\\",2):f(\\\"\\\"{8w@a\\\"\\\",2):f(\\\"\\\"{fJp*BKBGa<Cp@3bmbP.ipQtM<cCibRa20CclbSh+7<a\\\"\\\",2):f(\\\"\\\"},/beb:ncby,M<Sa|bd/Na+eU0A,Raeb+wXap|Va:o<aEa9b6b?aK/\\\"\\\",2):f(\\\"\\\"}bfbQaw;>a->8bj6F\\\"\\\",2):f(\\\"\\\"{.bQabqeuBav*Sai9FaV,6bA\\\"\\\",2):f(\\\"\\\"{CBN..@\\\"\\\",2):f(\\\"\\\"{u,u\\\"\\\",2):f(\\\"\\\"}3O?v>7wRa/1grwblbk*yb;0jrkgUu1bWaCcj+.|<aCr1o/bwb8\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{b:zzb>aOa2bRaabdopsFa2bdbkb>aRa=:T\\\"\\\",2):f(\\\"\\\"{*b?aC3Kscb/ujb?9P.Hs9bM\\\"\\\",2):f(\\\"\\\"}Uqcb+gOuu\\\"\\\",2):f(\\\"\\\"{fr=aubI.u3:|1bUaz4V*ShKv69S=1*Tsthh>E6-b-b+bTaph<a5;OnS29uM>e17bebL*-bvxt|:yC>Uufrlu*9y|M|Faz-j:=85\\\"\\\",2):f(\\\"\\\"}gu0b3b7353X?4u\\\"\\\",2):f(\\\"\\\"}8X;vyU\\\"\\\",2):f(\\\"\\\"}esBr?al7-b,5-0Mr3>dsWa407bm7a9fv9pvb;gTa+,55I1*3ipibJ8zb7=jozb3bjbs-1;GrM*Fa+"));
$write("%s",("=4q7b,8<8d1|bOav6\\\"\\\",2):f(\\\"\\\"}bG>cpapdw2xvfU+C*Kr2q<3uw,?j1Ba=-;-*pabh,tvo3Ta1bq7Y<DaAt\\\"\\\",2):f(\\\"\\\"}-./MribabhzB=Wamsgwwb>a>sAa2bEaCadpjofiE;UzCuT=hiB;D;r.ab<aK*23DtS\\\"\\\",2):f(\\\"\\\"}|bdbe=b.*gb.Xa6bwbssI\\\"\\\",2):f(\\\"\\\"}jk\\\"\\\",2):f(\\\"\\\"}blblr.qEa\\\"\\\",2):f(\\\"\\\"}wg4Xa|bDaBa*bfb8\\\"\\\",2):f(\\\"\\\"{bbdtk8ybWaB>ec5:\\\"\\\",2):f(\\\"\\\"}bC=Zai9ubQ5/|.b\\\"\\\",2):f(\\\"\\\"{io9k133X3K\\\"\\\",2):f(\\\"\\\"{CxEf4.*b/bR39bZambybkb\\\"\\\",2):f(\\\"\\\"}t4bN+K\\\"\\\",2):f(\\\"\\\"}2|dsd;4wibTa1p=aU-Ua8-cr=al7ibWa-bhbfbu/mbCap|dbf*n-y,9=c,f|Ty,x1bT*cbOn,rkuJxS\\\"\\\",2):f(\\\"\\\"{u/j\\\"\\\",2):f(\\\"\\\"}Iu7b6\\\"\\\",2):f(\\\"\\\"{*b@aw6<aYod\\\"\\\",2):f(\\\"\\\"}>ap\\\"\\\",2):f(\\\"\\\"}cbx-OaT1fbOan\\\"\\\",2):f(\\\"\\\"{-bqxDa-bGa*ycbkbL1h=vr?w>t74I-\\\"\\\",2):f(\\\"\\\"{*0b6b-bQa4b@a@yLgEaPa/|v*4bDrBuG+c3hia3693oQaxbjbQ1p8Na-bOk3b\\\"\\\",2):f(\\\"\\\"}bZ*"));
$write("%s",("ebg,74+bNav*cx2bPae+i,Va0bub:1/bubFav,hb>sixNw>a5;5b/b1bFaI-Cr6bNa*<A.o=\\\"\\\",2):f(\\\"\\\"{bzzv6DaCr5bzzPa3b@av*N59<=\\\"\\\",2):f(\\\"\\\"}Pf,b/\\\"\\\",2):f(\\\"\\\"{/bo*e53b3r\\\"\\\",2):f(\\\"\\\"{babtb8bNi3\\\"\\\",2):f(\\\"\\\"}dptbIwabXaRv-dabQ-;8*bGtJu=3k|FtybOaFt*bebd|atwb=/1bK7bbOaStcbh<lbP/@8Bakb;hd*dby\\\"\\\",2):f(\\\"\\\"{hb3oQ-4b,:\\\"\\\",2):f(\\\"\\\"{t8xe0H9w63o@wesg.*b-bYawbPxEa0bW7L,YaWa.b\\\"\\\",2):f(\\\"\\\"}/M,9bAq+bT9;87b|bH9i9u:xbxbYaUa3;CatbhbK7fb3bd\\\"\\\",2):f(\\\"\\\"},;\\\"\\\",2):f(\\\"\\\"}lw.39/7d3z\\\"\\\",2):f(\\\"\\\"}u.xxGy3bg.Tayb4bGy=aabubY-ubV:+2Ta3bSa@.4bjbk/=aWaPacbG6Y:jkRaFy+25b2br9xbBac1xb*bBp6\\\"\\\",2):f(\\\"\\\"{@aE6Ea/bWacbxbpq8bO:>a3bX,*319Xv9tmxA|Pw,5.hu/Eqgb\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}m\\\"\\\",2):f(\\\"\\\"}owT94b4b3j8b?acw>:e:;6wbDnAatbv/x,ivV,\\\"\\\",2):f(\\\"\\\"}bR1=adb\\\"\\\",2):f(\\\"\\\"}bT\\\"\\\",2):f(\\\"\\\""));
$write("%s",("}wpy8Xalb\\\"\\\",2):f(\\\"\\\"{bTa.b,bjbUqj*a4tpczWajblbitN8fb4b6|wb6buoib2yhbEacwubAahx8x5byu:95+\\\"\\\",2):f(\\\"\\\"}0c|QaYa8.U+vsbpF0Cx6-4\\\"\\\",2):f(\\\"\\\"}voRaXaubx3cbFa99wbws3oY7kb\\\"\\\",2):f(\\\"\\\"{9tqebibu1Vakb4a07Z2VzX2E+xb=v3oLgr8p8Fy?3lbCtbbn5jvmbus|*W/*b1,Ra4b:72jM4lbJ,cwd/WaZ\\\"\\\",2):f(\\\"\\\"{7bPaRavbvbmbdpl*T\\\"\\\",2):f(\\\"\\\"{g6\\\"\\\",2):f(\\\"\\\"{bl.=*<pecO|i*3u6bjoY\\\"\\\",2):f(\\\"\\\"{yyY\\\"\\\",2):f(\\\"\\\"{5bb+>aYaVo;qc|3ot1G6fbC3Dafb1bmbj5Pxlb|*zz\\\"\\\",2):f(\\\"\\\"}bqu>aY/zbm13oDaMv<aE.4bXaXaX\\\"\\\",2):f(\\\"\\\"{9b-bT\\\"\\\",2):f(\\\"\\\"}e\\\"\\\",2):f(\\\"\\\"}nvHvCo|gWa8bZabbz/c\\\"\\\",2):f(\\\"\\\"}N*cb<hUsLgUq2z5x,b,uQywsOy\\\"\\\",2):f(\\\"\\\"{bEaFaauZpJ3Gr,b0bYa024*u*M\\\"\\\",2):f(\\\"\\\"}kbkbW|\\\"\\\",2):f(\\\"\\\"}6X.h^127^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^32^[2fha\\\"\\\",2"));
$write("%s",("):f(\\\"\\\"})3(f\\\"\\\",2):f(\\\"\\\"{#v3rga(f;)0,73-c1bNv?7u3?7LuzbgbOk>|Cv0z=apqvbDaybYa8bDcxbhi.7Rrr5Lx3oFakbVyY/kb0v/tebRamh/bVaEad7.b*pZqGmWaTaGr@aSa8ba4e/SaVaSa?aN6RaL6db2bn-@a663oz-y2Ca7by2=6yyPa7b;6UambY\\\"\\\",2):f(\\\"\\\"{EaSa,5Pa>q:6Aae.EaqsTaVad4i4mbVa1bkpip\\\"\\\",2):f(\\\"\\\"{blbub4wkb+qmrZadb3/Jxlbiq|1XaOa*bGaW-,x-.jbwb/q@\\\"\\\",2):f(\\\"\\\"}Bahb>yRaCteu+,Oactx5C-<aezO5\\\"\\\",2):f(\\\"\\\"{5DambAacb|*3b8\\\"\\\",2):f(\\\"\\\"{8byoJu\\\"\\\",2):f(\\\"\\\"{bk0DaNalbe+6y:|-bkb5b91y*Qazb9b2b=a2byy3-St0wL4ub3bI/1yyymbztzb\\\"\\\",2):f(\\\"\\\"}b:|gbxtebabjtfb<y3i?aEa\\\"\\\",2):f(\\\"\\\"{bdpr|\\\"\\\",2):f(\\\"\\\"}lp5w\\\"\\\",2):f(\\\"\\\"}?0TpabEwNa=nfbN4XnmxXnRaibvqUaCvZu-.AnPt|0rs/bxbgb=vC\\\"\\\",2):f(\\\"\\\"{brAaBavbljjo6blbRaZ\\\"\\\",2):f(\\\"\\\"}Guxp*baxWayb-b|*ubOaSh<lVa?aOa<,NaybZa9te.-bSvvbBp3bhb-b6*ltdb7b;1z.vp3o-0tb3o\\\"\\\","));
$write("%s",("2):f(\\\"\\\"{tytz-xbMt4bwblrSa@aubI\\\"\\\",2):f(\\\"\\\"}m33bVa0rWalb,||bHnbbcoFa8\\\"\\\",2):f(\\\"\\\"}UagpQaR2G*=aB1ixf|Yai\\\"\\\",2):f(\\\"\\\"}d/Pavsc\\\"\\\",2):f(\\\"\\\"}QaibKu<\\\"\\\",2):f(\\\"\\\"}/sVa2qjb2b-pCt0bsygs\\\"\\\",2):f(\\\"\\\"}bRgZaQaicf\\\"\\\",2):f(\\\"\\\"}O0SaGr>r|b8b\\\"\\\",2):f(\\\"\\\"{bmbx\\\"\\\",2):f(\\\"\\\"{,rh/7|:\\\"\\\",2):f(\\\"\\\"}ablbjbszW|*bxsFthbXa5bcbqjbo/b+bipnh\\\"\\\",2):f(\\\"\\\"}lv\\\"\\\",2):f(\\\"\\\"}v.fix\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}lEuA0uc-b:.CaGa<.Za?a7bybvbYa:\\\"\\\",2):f(\\\"\\\"{lbibZa+bg,3oVs9b6222abq*h-+bjbOa0bRa9bFaptgbZazbNa@y.b\\\"\\\",2):f(\\\"\\\"}bjbL1xpgbr\\\"\\\",2):f(\\\"\\\"}1bm/mblbVaVaOaGtYaT\\\"\\\",2):f(\\\"\\\"}Grj1Vap0n0.bd1b/>a\\\"\\\",2):f(\\\"\\\"{*8bc*AafbPahbj|YaJ1,kc\\\"\\\",2):f(\\\"\\\"{6,El81+bRa\\\"\\\",2):f(\\\"\\\"}bOa-boh,-9\\\"\\\",2):f(\\\"\\\"{Oa,boh<jNaHzHtao4pFadb\\\"\\\",2):f(\\\"\\\"{bRaz/6-2p/1wbabwb\\\"\\\",2):f(\\\"\\\"{bxo@-"));
$write("%s",("TaPawbk|0bQm3zzb?o1rHzuw?af*ibxbT\\\"\\\",2):f(\\\"\\\"{Ra@atqDaCaebfb0bs-8bO.<jRa\\\"\\\",2):f(\\\"\\\"}u7b8bp,.hZpQa3babFayuSalpZaHzb\\\"\\\",2):f(\\\"\\\"{aoyb5zUafbjbxbcbR*CawbZao0m0Q*mb4b,x2b\\\"\\\",2):f(\\\"\\\"}lPrTzH+s.RavyJp>a++Ea@aFaP\\\"\\\",2):f(\\\"\\\"}PufbtbTaVoTaX*gb8blb//i04bvbf0d0Zp\\\"\\\",2):f(\\\"\\\"}bib\\\"\\\",2):f(\\\"\\\"{b+-mo|biqp\\\"\\\",2):f(\\\"\\\"}5bhbdbhc3bkb./-tDfybcbtbAa*uxt\\\"\\\",2):f(\\\"\\\"}bdbjbmbes4b7\\\"\\\",2):f(\\\"\\\"}xbkp,bk\\\"\\\",2):f(\\\"\\\"}-oZ+9bEaVaArXaTa@nwwVa2|ZalbAalbuydbXaabjbibebapEaAzb\\\"\\\",2):f(\\\"\\\"{3o*,OaCtAtox\\\"\\\",2):f(\\\"\\\"}bmb.bYa.bibPad/Zsab++In\\\"\\\",2):f(\\\"\\\"}w1bwbyb8b9bp,XxmbSaPagwAa/bjbgbf.gqWa|bxo.b2-3uyo3o5bOxCalb|bkbzb7blbYambehub2b|b,b<pub|bX\\\"\\\",2):f(\\\"\\\"{Stl*lbxbwprvSh8s4bRaww|b9+<aabeb|bXa\\\"\\\",2):f(\\\"\\\"}zJxkp-b?a8bydPaQ|ab5bbb=rBu\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"}UrBuS"));
$write("%s",("zI+zbdt@ze\\\"\\\",2):f(\\\"\\\"}=aUn,wtz@aWa=aSa.bRacb+bQaQa0-3bSh|-qpebjb5b-,Ta*b0zR+=am+-tF,dbWaC*D,\\\"\\\",2):f(\\\"\\\"}bA,eb4,?albnvbb.bWap,8bmb8bK\\\"\\\",2):f(\\\"\\\"}wb?a|gibCal,@aabHvnx?aK\\\"\\\",2):f(\\\"\\\"{/b3oNaOaAatxTaL*Ca?wubeb;j;xdbub3ok-1beb\\\"\\\",2):f(\\\"\\\"}b6bjbPa*bSaCa2r+b<a|gS,PaBqBaXzibubwoTuFaEaWawbPazbOa1btb2b+bkbQa9b@aEaZ\\\"\\\",2):f(\\\"\\\"}8pBr*bcdvuJz?n-tn,>a2rxwa,=aYafb.bKwh,0vabmbib0bybzbmbYa\\\"\\\",2):f(\\\"\\\"{bNaubVaCs*bXacb2b7bFn8b6bUagbQaBaEaNa|b@axhmbub-tO\\\"\\\",2):f(\\\"\\\"}cu<nVaFr/bBafb*rP\\\"\\\",2):f(\\\"\\\"}3bybabVm4aF+@uWru\\\"\\\",2):f(\\\"\\\"}kb6bHu8xSxZaR*4|AajkzpwbUaA\\\"\\\",2):f(\\\"\\\"{hbVvvbrhQank|rkbT*ioUgBv3byuvvBaShxyibgb\\\"\\\",2):f(\\\"\\\"{bzpSajzWaUaR**bVa4b*bib/tWaCa8x/b.bwbBzSqYa6bDaZu4b:\\\"\\\",2):f(\\\"\\\"}ubWatbluabgbbb+e,bPadbZaPaZzz\\\"\\\",2):f(\\\"\\\"{ebbb7bWa,bTadt-\\\"\\\",2):f"));
$write("%s",("(\\\"\\\"{sq*bjb*sdby*+b*b;z?a*bTawv<a?a3o0b*b>awvRa\\\"\\\",2):f(\\\"\\\"{*yukbNaY\\\"\\\",2):f(\\\"\\\"}Pa1bmqNa5bMvax@aXaaj;u8b7u5btbwb-p1\\\"\\\",2):f(\\\"\\\"}wbwbOaOaRawbebzbAyHzD\\\"\\\",2):f(\\\"\\\"}qvSa3bZaGyDawbbb3b,bub\\\"\\\",2):f(\\\"\\\"}b-o\\\"\\\",2):f(\\\"\\\"{bwb+vIqZa1b8b/q4bp\\\"\\\",2):f(\\\"\\\"{jb4bZa3b0vDavb<aYa\\\"\\\",2):f(\\\"\\\"}b.pf|ubc\\\"\\\",2):f(\\\"\\\"}7bCrSa1bSa7bgbcsebPoRzzx*lAuBuenQzjx+bybUaZaeb@a+bwbcblr9b\\\"\\\",2):f(\\\"\\\"}bkbe|ubXaebwbkbCsgb:\\\"\\\",2):f(\\\"\\\"{YaNa\\\"\\\",2):f(\\\"\\\"{b6bvbjoPaXa\\\"\\\",2):f(\\\"\\\"}bYa|bQnvbJnFaxs-bZaewZp*bwy3ot|mbtbtu,bOalbkbpoUa3obbZahcTa\\\"\\\",2):f(\\\"\\\"{bqjlb4b5t\\\\\\\"\\\"),\\\\n(\\\\\\\"\\\"Qa\\\"\\\",2):f(\\\"\\\"}|\\\"\\\",2):f(\\\"\\\"}w|iCa|wvbbbab=v,xFaOa/bcbhc>aDp0pXa;q,x*buzebtbeb4bxb=aybKxlbWaabwwdbJxvbOafl*b7b6wBq*b/gSaKx*b,uCvEa+b5bwbFaXaIw+ibr6\\\"\\\",2):f(\\\"\\\"{5b*b2b1babvbVahw+\\\"\\\",2):f(\\\""));
$write("%s",("\\\"{GzEzCzAzbbDaUaSvQvc\\\"\\\",2):f(\\\"\\\"{nvZz0bXzSaFa.wOzNa\\\"\\\",2):f(\\\"\\\"}zcrzzxz|bjkYakuZpmb;uabEaeuwb>pHz8b7bes.oCt\\\"\\\",2):f(\\\"\\\"{bBu*xSoyx|x\\\"\\\",2):f(\\\"\\\"}l\\\"\\\",2):f(\\\"\\\"}xwb=a:z8z6z4zbb,k\\\"\\\",2):f(\\\"\\\"}b-bTaUg\\\"\\\",2):f(\\\"\\\"}bWaYadblbfpIhlb>aNa.b1b,xxbhb,bFavblbic*bOaazlb0wNa6b4bYa*ttbtbBa\\\"\\\",2):f(\\\"\\\"{b+bcbAavbiytbmb<aFaDvky4bhbYaOt4y2y0bAaabYabbVa\\\"\\\",2):f(\\\"\\\"}bPa2bCa:pwbXaRa8b>p|bAa7uDa1y;pbyVa8bwbUptbUaauUaOaky|biygymbgb4buvzbkbAa.bDa8b4bff|bwyuysyShHqeb0wVxyb3oDp|bgbib3bCa3o2bAa,p=aOajb\\\"\\\",2):f(\\\"\\\"}bdviu/bAaWaMwKw4w/vcvkbBaWakb2b5b8x*bQaabib.btbmtWa1bcb3bjkbbcb<a1bVa6bYa,sPw,x7x?w-b@wab\\\"\\\",2):f(\\\"\\\"}bNaYaZanvdjZaCa,xhbBatbgbPo\\\"\\\",2):f(\\\"\\\"{x>uZmBuDuTrUm7bXaPaTqjbNa\\\"\\\",2):f(\\\"\\\"}b5oPaub7bjtkbmb0beb.bjkShXw6b+q5bdbMr*bRatb?a6b8b-t8bAaXaAa\\\"\\\",2):"));
$write("%s",("f(\\\"\\\"}b3bYacb/bdrgcdugb\\\"\\\",2):f(\\\"\\\"}bDrSh:w-b3o\\\"\\\",2):f(\\\"\\\"}b2b,b3o.rrs+b6bZafbUa?a1b*qSaZpubbpmb5b@tdb=a9pabhsCa4b8b+bLgow,pdq*uWa\\\"\\\",2):f(\\\"\\\"{vgbYoPa9bbbwbgbOubb0bwb8bcbCawrmbjbdbzqUs0b.b<ambxbib>a3o|b-snr|b4uybkoQa0b=aebFaZl2p5bNaXabr0pEaetBabr\\\"\\\",2):f(\\\"\\\"{bUaPnVsYatb7uUuNatb<q=ogbeb/bmbNazblb0bXa-b/bkbabUuBagbqj1bfb\\\"\\\",2):f(\\\"\\\"}b0b0b@a|bVatbfbwbWa*bdbxd2p7b.bBaZi6tcb6bmgIoibbb5b.bOaXaBu?uNoWmVrSrPoToOrqqAajbShoq\\\"\\\",2):f(\\\"\\\"{b/bsq*ueb5bEaubysEs*bEaYa0bkbOarp/becZawbJd=a*b+behKtOacb1b7bdj8bebXaDa9htbgcSaubxb7bZa.blb=acbCtZa2pab2b8bipxb2jSaUatb8p8b/bXaZahq0bcb,b=aCa-b@a*sPaArkbFa?a/b-bRaUaxbEaooQpzbcqdbmbQalb3o\\\"\\\",2):f(\\\"\\\"{bWaXaNiOauo1bXpQa?assBsAadbgb,b6bTaab4bbs=atbNa3b5byb@aBaxb\\\"\\\",2):f(\\\"\\\"}bzbTaFa7bir=pWa3b,d@r2b.rubfbErtb@axsvsGr\\\"\\"));
$write("%s",("\",2):f(\\\"\\\"{b4b6bFaYaeb.s4bPaNa3o/bPa.bbb,bqrDa@axb.b=a8bdber3bQa7bWq@a8b.bTaQaSa\\\"\\\",2):f(\\\"\\\"{b?aab^127^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^32^[2fha\\\"\\\",2):f(\\\"\\\"})3(f\\\"\\\",2):f(\\\"\\\"{#v3rga(f;)0,73-G~Va-bfoUaXa9bqr2jVaUaTaBacbmbmbXafbvb0bVmhiQrcnPoanfihiOoRo0b3o.bXaUabdkombzb@a-bfb|b6b>abcmbUqTaRabb:nzb?a\\\"\\\",2):f(\\\"\\\"{bEf>aebvbTaCabc\\\"\\\",2):f(\\\"\\\"{b1bkb9b.b?aebTa2bUaGa?qRaBa.bAoTnybmjdbcbWa0bFaSakbTalb5bOaubQa\\\"\\\",2):f(\\\"\\\"{b.bUaSaRaubjbcb9bzbjbRazb2b@a2beb;qAn3olb@aEq9bfb-b3bUaSh2oVazq7b2btqrqpqXa.bkbUavb@a?pvbZa\\\"\\\",2):f(\\\"\\\"}bRpiqdbwb\\\"\\\",2):f(\\\"\\\"}bDotb4b,b7b7bdb0bPa,babxb3o,blbUaQa>aib,bebVajbjb7b0bWaBaFaBoab7bUabb\\\"\\\",2):f(\\\"\\\"}bebmb3bmp\\\"\\\",2):f(\\\"\\\"{pypzb=auphb*bBambPa|bEajbFaPaCambFa>aTafbibOaCajb"));
$write("%s",("hb@aibkbcbibjbVo7btbbb|b2bEo|bmbBaDakb=ajbyb|bSaZaFaDa4bDaFa.bAa0bZaDajbTa8bOaTabb8b5bebhbcbwbVmPo,lMoIbfnYm:ibnebDaEl6b6bebDfkbdb+bSabb>awb*bCa<a|b<aNagbvbNa1bGaso7b<a>aWnSaXaFagbzo\\\"\\\",2):f(\\\"\\\"{oyowo/bYagb7bAaFaShqbjb>a=aAnCaxb+dXabbjbpmnkEaao/bUa>aFaVa6hdb/b2jeblbzb,bNa7bvbCaEahb<aCabb*byhQaub*bWaQagbSa,bEa7b6bAaEaHl,nSlsnlnjn>fzmqm6g\\\"\\\",2):f(\\\"\\\"{n;asnrmpmjnrnDlwn2mSgwmKmwbic8aNm9m9lmnEaDl:mgm-a,mcmamhidn.lfiXmVm9aVmVm+l4a/l/b\\\"\\\",2):f(\\\"\\\"{f-a|hub.h|eEm=m0mAm7l9aEaOa1lim:lwmIlmm=g:a2m=aAawm/mCaSljmum@a<a-bzm*mJlzmLl8lvmymAa:aCa8asm>aKlClRlMl>lUlAa?a>aJl|edmzb;lOl<lFlBa8lBl@l*bvbtb/b-aJdHd1lNlElJlHlSe|eAlGl?aAa-a7l8a=l;lFa@a8l\\\"\\\",2):f(\\\"\\\"{b6lHa4l9a|e5lxb8a+e-a1bDf1lrl8arb8a>fhi-lfi\\\"\\\",2):f(\\\"\\\"}l3a9i\\\"\\\",2):f(\\\"\\\"}lgikl<h<g6b-a+czbxbubHaqb6aqb2i3"));
$write("%s",("i1i5aqbvg-aff1bzb.b;gnbxbjiShDgBgUk@jobjhwhbkwjZj?a=a9isi2kxi0kbh.ktcBa8i|b|bvbAihc6fJjakFjBa?a8i6e|hrb3b\\\"\\\",2):f(\\\"\\\"}hKjTj=ikhGjDa?aDj2b3b4i;f+c/g-a=g-b0jCa3aKa\\\"\\\",2):f(\\\"\\\"{b;aigwbccIa3b1bmj,b|b0abhxhbhyjRjujCa8i.bbixh2hIj<i:i@a8iyb3bBj?a>ixjuivjBa>a8iPcri?j1aHgsbubwbSh-a1j/j:a;b,j1b0b-b3aAa3a7b-aSh.a:b:b,bxhkhwiPaUh;i@a3a|hwb+b-aPcaj/b8b1bPcxb;a;f-b0gZaNf|b.b5b-aSi+i3b=fvb|b+g4iNfEf3bgf;a<b:b3b-a8b+g,bxb2b2btb;axhEhviEh3a>a3a5anb-a2i/b3b4b.bHa8byb2bhgtb=fxb5b+bCgxhvhThGhvhGg=g;gHaniniFaGaRh|fld4a/aei-f4a-aEfCfMaFa=aEh-bGh2h1hGa+bJd?h9a/b5a|fCcng-bPaBaob2h6aKaMa9aMaIa5axb3b.b4b0bxb*htbDfxhHgvhGaMb*g2bzb;azb-b<gccJa7b?a?aahkhCdYaOaVafbVaibNa=abhbh?a;a6gVaNaUa/aHgahHgvbpbEa*c7b@a>aCaCa>anbJdubSczb6fMa-fob,fyfwfuf2bsf/a?g-f;d+c1b/bNd3bHa?e-a/a,f:aIa+ctb"));
$write("%s",(",b:avbldub4bcb-biggcfgHaebdbJaGagfef8a1bxbwbtbxbUaac|b3bCffb-f-atbxc8f?a1a-a6a5bGf>azd:a,cNaGfwb.b;b>a1a,c:a-a.b\\\"\\\",2):f(\\\"\\\"{bvbxb5a1a5aCe2b-a:b1dtbHa6a/c2b3dMd-aDdBd@dmf/aob5a.d,d*d-b4b7eSc;axb+b.bbcZb0cbfJasdHa/aed+e0cGb/d,btb-b4aWbudpcgdLc=chchd6areOapc0cNb/a;bje/eGaHb5dedOb.a8aNd8aLdLa=a>aIaOaJapb6a+e5azb+cdcfbhc;aOaFdYd6aHaCa@aIaQd8aHa=a.cIbCbMd\\\"\\\",2):f(\\\"\\\"{cycvcocRapcXbocTa;b;bpbgbYdJaGbRanbQaJagbnbcb>dqc5dpbebnbOa8a0c4aJaTa5a+btb5bxbJaQa,c*cRa5a1bzc6aedMa0c3bldjd;aeded8ard5a6a5aedxb/btbvb2bxb,c1b4b3bxb1b0cocPa8aNapcMagdUc3b|b+b/b2b4arcFbnc4a=a?axbtc4aSbJcPbKckcic+bZb3b-bzcXbqcFb5aMa/ancvc+b+b|byb4a9cVbNa5aRb7cFbnbFbMapb2c.aMaFb.a4a5aJaOa-a-b|b-aeb5aicybHa<b/akc>a>aXb6aOb/a8a6a/apb4a1b.b3bvb4b1b3b2b-b.bvb4anb/aJaPa5a8a4a6apbEb5a5aBb,b9a4apbpbnb8"));
$write("%s",("anb4aGa=a:bJacb!PQ1ca61QQ.ba~[2xha=s,y=z,54[54%.4[e6&yay,]99999[gnirtS wen=][c n3aea\\\"\\\",2):f(\\\"\\\"{)v]y3b&a(niam diov citats cilbup\\\"\\\",2):f(\\\"\\\"{RQ ssalc~5[~5qfa cdlnl3c/a;maertStnirP/oi/avajL tuo/metsyS/gnal/avajq5bdateg@3doa2 kcats timil.v3dga]; V);U5aC3ecaL[f6aa6hha dohtem?3e;4nga repus&3ecaRQ@3cgassalc.@6[@6ioa(=:s;0=:c=:i;)$5ajaerudecorp34[34eqa(tnirp.biL.oken\\\"\\\",2):f(\\\"\\\"{24bianoitcnufc:[83\\\"\\\",2):f(\\\"\\\"{martStup=niam^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'>3(ba7U3vJ4vba7I4.da,43?4[fa(f;)5/6/#6[#6[#6[#6moa(etirw.z;)tuo.-@aba(q?b~auptuOPIZG.piz.litu.avaj wen=z|5[a7["));
$write("%s",("a7;ca94A4.l41ba0j4[w5ada283m4[x5[x5[x5[x5[x5[j4(da373x5/fa wohsP=[5?[5?;ba35?[A8[Z:[x5[j4vea1982m4.batv9[V:[?4:da12927[=8[V:[x5[x5vca04V:/5aR0Z0Z/512152353/2/2166263=4/3141726??:1518191:1/I9[.;[?4:da063eT/r9[/;[x5[j4Fda66957/da*6 .C[Z:[?4;da348Z:[A8[Z:[x5[57wca8457/ea1312aC[a;[?4<da423VF/C8[a;[x5[j4Fda200a;/YB[W:[YJ<ba1OV0>8[W:[x5[YJGca15XB/fa41310\\\"\\\",2):f(\\\"\\\"{9[[:[.[;ca92B8[B8[[:[x5[x5wv5/qa;t:\\\"\\\",2):f(\\\"\\\"}%%%%\\\"\\\",2):f(\\\"\\\"}fi\\\"\\\",2):f(\\\"\\\"}*-84OH2ca7786[86[Q8[x5[QPwba9R@/(a]i[\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"}+17\\\"\\\",2):f(\\\"\\\"{<84.;i:-i602\\\"\\\",2):f(\\\"\\\"{;i:911\\\"\\\",2):f(\\\"\\\"{;j:6323?[tA[?4:da550d9/xa(tnirP.tmf\\\"\\\",2):f(\\\"\\\"{)(niam cnuf;V4[;6[;6;ba93;[><[j4gca69mO/datmfY6[>8[5R;ca5847[?8[V:gca02?80saropmi;niam egakcapo7[O8[?4;L[1ga(tnirp[A[+6[?4;ca36(I/|"));
$write("%s",("<[j47da444l4.ba-W6[<8[i<[A?njanirp tesnw41ca21T9/la1 etalpmet.f6[F7[)L<l;/ga(ntnir|D[*6[?4;ca93SG/baf)6[)6[?4?ca11EG0$a,s(llAetirW;)(resUtxeTtuptuO=:sc5[C6[?4;8=/#BaC4[(6[(6[v3kdaS C&6[&6[*D<3=/ca&(?4[$6[G9[v3kba r=[)6[)6[r=[&6[r=[83)iaRQ margoP9[-6[-6[P9phaD : ; RW9[-6[-6[v3mba^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'>4[#6[#6[#6[#6[#6[#6\\\"\\\",2):f(\\\"\\\"}i=[$6[$6[v3lqa. EPYT B C : ; A36[36[36[y=[#6[#6[#6[#6[?4[#63ka)*,*(ETIRWs=[.6[.6[G@nhaA B : ;,6[,6[,6[v3lba [2cF4[+6[+6[T9oia: ^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\""));
$write("%s",("\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"' ohceI4[.6[?4[73kpastup\\\"\\\",2):f(\\\"\\\"{)(niam tniL4[164ca01?4[?43ea%%%%@4[%6[?4[%6[%6[?4[73\\\"\\\",2):f(\\\"\\\"}paparwyyon noitpo26[M45<4[<4[<4[<4[jD@hanftnirpD4[fa(f;)3D4/kaetirwf:oinu41ba2u4.ja>-)_(niamt4[Q8[<4fWP0gacnirp(C4-ia(stup.OIK4/rKajaM diov\\\"\\\",2):f(\\\"\\\"};)B3(ca11g62oatnirP)--n;n;)sn3a<a(rof\\\"\\\",2):f(\\\"\\\"{)n tni,s tsnoc gnirtS(f diov\\\"\\\",2):f(\\\"\\\"{noitacilppA:RQ ssalc[k4rga@(tnir>MblaM dohtem06x*3cl;abNcuadiov;oidts.dts tropmtNnra1(f\\\"\\\",2):f(\\\"\\\"{#(rtStup=niam&3kkaenil-etirwb8dva(,^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\"));
$write("%s",("\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'s%^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'(gol.elosnoc;)^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'73g\\\"\\\",2):f(\\\"\\\"}a^129^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):"));
$write("%s",("f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"' nioj.)1+n(yarrA>-)n(=fI3cva^31^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",2):f(\\\"\\\"}54,1\\\"\\\",2):f(\\\"\\\"{.^127^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"# qes-er(K7c.4cba^31^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"p3lg3fw3hla1% ecalper.j4dea^128^gXc/arts(# pam(]YALPSID^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^127^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\".NOISIVID ERUDECORPA3cma"));
$write("%s",(".RQ .DI-MARGv3g53d|bNOITACIFITNEDI^127^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"[tac-yzal(s[qesod(^63^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"))System.Console.Write($^63^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"Put caffeine \\\"\\\",2):f(\\\"\\\"{(int)c\\\"\\\",2):f(\\\"\\\"} into the mixing bowl.^64^n^63^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");M3pva^63^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"Liquify contents ofE3oeaPour^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",72):f(\\\"\\\"\\\\"));
$write("%s",("\\\"\\\"),\\\\n(\\\\\\\"\\\"\\\"\\\",49):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'3w^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'4e\\\"\\\",2):f(\\\"\\\"{abaking dish.^64^n^64^nServes 164cma\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}^31^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");\\\"\\\",2):f(\\\"\\\"}/****/e3a^15^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"),s[999999],*q=s;int main()\\\"\\\",2):f(\\\"\\\"{int n,m;for(;*p;)\\\"\\\",2):f(\\\"\\\"{n=(*p-5)%92+(p[1]-5)%92*87;p+=2;if(n>3999)for(m=(*p++-5)%92+6;m-"));
$write("%s",("-;q++)*q=q[4000-n];else for(;n--;)*q++=*p++;\\\"\\\",2):f(\\\"\\\"}puts(s);return 0;\\\"\\\",2):f(\\\"\\\"}^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"))\\\"\\\",2):f(\\\"\\\"{s+=^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"00g,^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";for(m=1;m<256;m*=2)s+=^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"00g,4,:^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"+(c/m%2>0?^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"4+^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\":^7^\\\""));
$write("%s",("\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")+^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\",^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";f(s);s=^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"4,:,^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";\\\"\\\",2):f(\\\"\\\"}f(s+s);for(c:Base64.getDecoder().decode(^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"kaAREREX/I0ALn3n5ef6l/Pz8+fnz58/BOf5/7/hEX/OZzM5mCX/OczmZzBPn5+X/OczMznBL/nM5mZzBPu++fPPOc5zngnnO"));
$write("%s",("ZzOZgnBMGAW7A==^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"))\\\"\\\",2):f(\\\"\\\"{c=c<0?256+c:c;for(i=0;i++<3;c/=8)f(c%8);f(^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"8*+8*+,^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");\\\"\\\",2):f(\\\"\\\"}f(^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"@^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");^1^\\\"\\\",4):f(\\\"\\\"'|sed -e^1^\\\"\\\",4):f(\\\"\\\"'s/^16^/^32^/g^1^\\\"\\\",4):f(\\\"\\\"' -e^1^\\\"\\\",4):f(\\\"\\\"'s/^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"/^16^q/g^1^\\\"\\\",4):f(\\\"\\\"' -e^1^\\\"\\\",4):f(\\\"\\\"'s/"));
$write("%s",(".*/print ^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&^7^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^8^nquit/^1^\\\"\\\",4):f(\\\"\\\"'^3^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")\\\"\\\",2):f(\\\"\\\"}^1^\\\"\\\",121):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")\\\"\\\",4):f(\\\"\\\"');\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\").split(\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",128):f(\\\"\\\"^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");for(int i=1;i<a.length;a[0]+=a[i+1],i+=2)\\\"\\\",2):f(\\\"\\\"{a[0]+=\\\"\\\",57):f(\\\"\\\""));
$write("%s",("\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",185):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\".repeat(Integer.parseInt(a[i]));\\\"\\\",2):f(\\\"\\\"}System.out.print(a[0]);\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");\\\"\\\",2):f(\\\"\\\"}\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";FORiTO UPBtDO INTn:=ABSt[i];print(REPR(50+n%64)+c+REPR(50+n%8MOD8)+c+REPR(50+nMOD8)+b+\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"J\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"+a)OD\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans c 0\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"do\\\"\\"));
$write("%s",("\",2):f(\\\"\\\"{D(Integer(S:get c))\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 35 39\\\"\\\",2):f(\\\"\\\"}(<(c:++)(S:length))\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 24 149\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");end;\\\"\\\",1):f(\\\"\\\"\\\\\\\"\\\")\\\"\\\",1):f(\\\"\\\"nsys.exit 0'}\\\\\\\"\\\")\\\"\\\",0)]]></xsl:template></xsl:stylesheet>\\\":s=\\\"   \\\":For i=0To 7:s &=Chr(32-(Asc(c)>>7-i And 1)*23):Next:System.Console.Write(s &n &Chr(9)&n &\\\"  \\\"):Next:System.Console.Write(n &n &n):End Sub:End Module\")\nput=s\nprint\nqa!"));
end endmodule