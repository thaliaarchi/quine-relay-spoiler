module QR;initial begin $write("%s",("Module QR:Sub Main():Dim s,n,i,c As Object:n=Chr(10):For Each c in\"<?xml version='1.0'?><?xml-stylesheet type='text/xsl'href='QR.xslt'?><xsl:stylesheet version='1.0' xmlns:xsl='http://www.w3.org/1999/XSL/Transform'><xsl:output method='text'/><xsl:template match='/'><![CDATA[write,format=\"\"%s%s%s\"\",\"& VbLf &\"(\"\"\\\\write{-}{txt}{(\\\"\"with Ada.Text_Io;procedure qr is begin Ada.Text_Io.Put_Line(\\\\\\\\\\\"\"print\\\\\\\\\\\"\"\\\\\\\\\\\"\"STRINGz:=REPR226+REPR153,a:=z+REPR166,b:=a+\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"2\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"+z+REPR160,c:=b+\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"8\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"+z+REPR165,t:=\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"write('implement main()=print(\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"BEGIN\\\\{s=(\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"#include<stdio.h>\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\nchar*p=(\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"Ra#include<iostream>!nint main()\\\\{std::cout<<(!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"class Program\\\\{public static void M83apbSystem.Console.Write(!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"let f(c :Int):Latin1=if c=127then!!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"!!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"else(string_of c@!!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\" g caffeine !!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"@$3kEa!!!!n!!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\")@f(c+1)in print(!!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"Quine Relay Coffee.!!!!n!!!!nIngredientsq3aha!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"@f 10U3cgaMethodz3c#a);let g(String ->[])!!!!n[c;t]->w4edaPutY4spa(int_of_char c)05auainto the mixing bowl|4ejag t!!!!n|_ k4gtaLiquify contents ofE3oeaPour\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'3w\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'4elabaking dishv6biaServes 164doain g(!!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\")))s!![2aca!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\" [2bo3cparts(nltnirp(])]v3cja.NUR POTSp3cx3dp3jba!!M3dp3df4fda[))j3ci3e,3cp3l[2kga\\\\};)06xu3kgaqp]\\\\}\\\\};@3\\\\}ga)1(f\\\\{#+3~ba3+3&ga7(f\\\\{#.,3~ba5&4\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'ga13(f\\\\{#+3O97l,3tkaD ; EYB RC73(da,43.3\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'daDNEZ3Sda. Ab5VeaPOTSc5Wb5TmaRQ margorp dS@aj4ObaSj5UV3Lca36V3Vba&P5MX3agaS POOLi;Vea\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'&,)i;Uga. TNUOf5Tfa(rahco7Nh5cgaB OD 0l;Uca&,t9Rca)At:Vo:UiaEUNITNOC0KiyIzga(tnirPLI(ca01q9Uj9Vm8OxCceaRC .b4Ska,1=I 01 OD3GWcaPUc4Tw<Rva;TIUQ;)s(maertSesolC;4Rmr4<la721(f\\\\{#n\\\\})8i3ag4Mda552X3Qia115("));
$write("%s",("f\\\\{#\\\\}Y3Mla3201(f\\\\{#mifS>$g7*da402h7cj3bh7Mpa904(f\\\\{#;)\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'\\\\})2392:\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'?A-da354w9aka\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\',\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'&\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'(rt.\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'%6Mda957v6\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'k5-ea7331RW,y7,eaq\\\\})6j3bh4TE@Oca51h7Tca561>aca\\\\}\\\\}2<Nb6Uj8[ga!!!!\\\\})19s;Uea5083h6Yea&dnek8[w?Iba3VH(w?.ca59l9[t;[$a\\\\{#&&&PUEVIGESAELPn&&&&1,TUODAERs3a$4Mca77<?Uea1232:>[-8[g5Oda745g7Tda945BVa$a&&(etirw;\\\\};u=:c;))652%%)u-c((||\\\\}6[)8Rca33d?Uda167*9[T>Uda#-<b5[FTG8S)-R/a4a7>[l8[ea&||iz=Nca78n;\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'=?.ba0q=aEC[m8Qda307FYVGZa\\\\{>YhaBUS1,ODv;[p8Qda2349SVca66iL\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'i6[q8.WHbma)3/4%%i(&&&&HT[KXHca70zPUea52034>[\\\\{OVba82>a=BRba1~9b0US(;[n8Xda7270?Uea96312>[/TdNa2=:/t;2%%t+2*u=:u\\\\{od7 ot0 yreve;i-=:u;1=:+i\\\\{od))1(evom(d"));
$write("%s",("ro=:t elihw?s;)s*jU[e9Tca51%?Uda149i9\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'i6[kU1IIPca19~@Vba5~@aw?[*D[ZPLba6v@Vca33v@aJJfi6[q8[h4Lba4%?Vda062\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'>[nb&n&&&&dohtem dne.n&&&&nrutern&&&&V);gnirtS/gnal/avajL(nltnirp/maertStnirP/oi/avaj lautrivekovnin&&&&u9[Y3Fca95+@Vba7~<a,?[t9[jb&&&&&\\\\}\\\\}\\\\}\\\\};0=q;)]q[c=z(tnirp.tuo.metsyS;)0(tArahc.y+z=]++n[c;y:]q[c?n<q=y\\\\{)0>2%%++i(fi;48%%)31-)i:3c&as(+87*q=q\\\\{);45951<i;(rof;n)rahc(+>8Mca71cBUda719lF[>9[AZQca59sJUba414a?:b[2cl6[t8Qda808OZVba86Q[T?Z[2coa=]n[c);621<n++K>aqa0=q,0=n,0=i tni;35[Y3Gca33R?Uda1677E[=8[=8mdd6a2b9anm2a4a5azb@d;axb,A2b-bt\\\\{Ga6aUcYfLa4aqc0cYjyb4aJaJaYf-ayb9C/bq5Hagdgdrf;fHawb;f6apb7b@lnbCbTf|bmn;dLb>aSi2a6a|bKaKa6abm:a@aEa2avb5a5aveHaAaGay>=aJabcXbVbjc+hDhzCCf3b8V.d>6JaMa\\\\}bJaPaCf@WJaJarcJaJaTaJa8bqo;a8"));
$write("%s",("bJ*Kaj.b1TaCfRrKUqOZ\\\\}Ka8bqO?aTaj.j.b1zCV\\\\}JaLaJaj.8bNaf4cca8b)9Qua(f\\\\{#NaeszC:b+b3b+bCfe3aka\\\\}bJaHaJa8b<4a+aHaJaJaQa?O;a8bBN:aUa:aqoCb2fbcZbXbVbwbk7gea>a8ao7aoajcms*bjc7aCbTfu7aoa+i2a6a\\\\}bKaKavbg7aVa=a*m:aXFJadczdUbCcohjc7aEaqbCcKgsbsb;dLbTb2fObldidpbjcHagdidpbrdCc8d=a-a<gbc3bJcrm3bea|b9ai3fEad7apb>yJdHdRihc1bZ1Jb|cV=Rhlx7a>y5a2bIgMa<gbc.dhYJa>a2a:b6a5a-bBy3biaGe/pvc6a53k&bJcMcvbvckd=a=addqelbOa-aRalbOar2UpteQdfeteGh7b3f|hMiHh*f.f;fGhGhUc>jFkKhg+-bjh9a4aSeqgig7hTh/bJc;a\\\\{eWgaj2f1b4b3bJcEgKg-eQ;c/a9aWhGh|k2a-ejpGhte>jwh4aMiHhdh4f*fZf7l0bMe\\\\{3c#aMf-h8d*fZfJcGhXgyeUcOkQhjb7emxk=ahbLN;a,bRh0\\\\{fbpbreub6cXblr,bnbreCep6,fCe.dhYzh-heh7hVhEaEdajAf?g=gHf9a7btcCeuI,b-b=g3a=a9a7bubxbu3g93gea3aAa;3kM3a93kha,b9a7bm+3fmacgCaBa+h9ae,/3ciag*7n3bVg73aca3bm3a1aCe+b"));
$write("%s",("Bd@d\\\\{e=g3asb>gAa3aMeGhXeqgQghgOgbg>gEa3as3gcang@6claSeqg,h;glfMaBMxa52(f\\\\{#(ntnirpn\\\\})821(f\\\\{#~>#n40dae=aO9gU5icaMgQ5inbvXGfGhlf7eGgZf9agxkP2a2a7uThkg1i.f;fMeGhu88aGhpbhgHh*f2fJaJaubve3fKgCe=anbre3flgyb6g-e,bJaGh7b5a*fZfI3cA3esa9a9b9aMg3flgCeGh>aq3aea@a@as3c-au8:a|b9a0b9au87aGhu8Ia|b-e:a9bJa0b3flgBjU3c%aMg9aCaAaJa9b3flgnbreJaEgoh-e,bMeo5g/a-ea:CeDdMfidpbreqmCeqmCeEggf-e7n+dCeqmnwbbw3aeaGh7bw3iqaqmnb*fDg\\\\{fZAJc6a04a4a8b9a7b-eMaJayb>a8qGa*mJa|bCezdMelfjfJa,bJe*mJa-u3b,aGhGhu8p,-e+b|bOc:a+hJaub-e.dOc?ag+-bJa30>jiashqh3a3bJ>ii;aoa*h3aBrGe=g*h3a>8eBj5h3h;awb;fGhqmv+-d<ioi4k/j2kv+MeciIi-k+kEkNkjiEkxivbm>D2tbk8gDQtG?Oz<yxVjbZaxVSw+ys1*.7?8BEaQu>aGT\\\\}oanHyEaB0gVuCBaEa+x2rMhwnqqIvA+Uka*Nl|W1bgbhb>lhb<abnhb>aEBP:xpYa|Wubhbbv8m@aXa+zZl.mR=gVa*RlLP6@:GdmP\\\\}Ba"));
$write("%s",("ibOKWqP6zt,bm,x+mb*t|b=aaNMqvp\\\\}rLNEa1lEaP5nESag9WlrwvXO\\\\}t1Xa75eyRv-\\\\}.6gQwnyxop0+/+AaxbC\\\\{B+tm/bRwpPZjgklP1Yj.bv-oLmuIYafl6b758b\\\\{tnBGvHEZ\\\\{ubhr*tq5+:yNXPR1clOK<sg*hHp:k4ZZwsDL,bbzrlabBX-\\\\}@sVpkbibO7Qq,\\\\{D2=DvbDa+wYlME9PxTVw:D;LgnPa2rYo0f/bjBxb|-Ynyb-*T-N-a;=a+9W4uufbOaoq5tu5EwvpCagbabNat;;qq5Gp-b8rkh>YKzEa5--d4RAaqWRIQIibws.oL:yXJo8bMu@8*bJokhBp/sCagbQu>aulJWxb*bXao\\\\{soSwLulqfT=wPawlDEa5p;fCvbv+DaZHplt4dt01L@\\\\{tJo\\\\{bqS,XSzm1Aw0lJQllAdIvA+R=qcd4A+Uk7v-bE=BaEaDlu2eD0ylbdl7N;LqlSarlplnl;OLy1=/=\\\\{m>aLv=a,bK:|=Gwi3mbhmsQo*zG>ax>iWEa,Xuben0wl=1b=2SNu*C-*t*b\\\\}pFw+;2BR=YaoJGmdlA?Za/bgA3bi=MZMp8mb.ibVa*tE-R+5Dib1EW3xb\\\\}BjluyBaEaw59slbl<blYlztGObl*bNl*be3aXbYlztvb:29o5>lb@aPa>y,Kg<Vd8Jv+J*2b<+Jo:MPaEaA:k<hlGdK;Ea:AFwHN5>lbE-Xnh<FartCafn+2O;klqsK;fn"));
$write("%s",("Zu\\\\}s\\\\{SLC75EaI-jlN@BaEa@aK;6XdbjlDlUa;;J*hriWEa\\\\}BjlF-R=\\\\{;UaLCQ;JsD*LC<a8bGnT\\\\{9We5e%cNabva*mbDa\\\\}>jlRmhm7biWEaRm5ndb?mZ:hbCaFx>uFxrwYa\\\\{s/=8xs-9WAaztMtcwgD\\\\}C.bIy9pem\\\\{.AMR*lv0@>:=a?vhb:5vbYOC8H\\\\{blm,pA.bdzL\\\\{|\\\\{mb,w/oLr+IIdDa?dYaOSmbCL50<aub1bhb6b=aDa\\\\}N@?-mX,o8F5ACk<-mX,hbNaCaI5V9u/qohbNadz0bN9DL#3c1fRanrib=a,b-b5m@9:ET><a9=9r3m+b>l<l?ajbZ9Hb50/=7cplrrB1jb?4,mQ9DaulA>jbGCYW?aafhbo9ql+rtrou1l\\\\{oQt3?H;nBabJmeXs\\\\{9bfvy7xlQahbPaU/Najb*t5+,G\\\\{subimU/C7ZvZvx0+0.thYfC?5hbSPGTj+R10wBmjB2mmNdx<tyN?.-bVUiy:X+XvXI5*CB6dzwbK;gklP5Jhbd-bbbStbx?2:cb4hB*zme*mbGdDa\\\\}0\\\\{sF*DaR=5/5/7eT8||a\\\\}gtrS:M\\\\{+t.\\\\{+|1wbGa*mzbVUT>RtUEYW?a5YD3J9?4|l5x7bCaub-zfWjI+UImrSUlSl*zD3HptG2QC/*0Aa8.mQ9E*b=aFaqAf6FW\\\\{RUl9oJ10.DHUagSJlg|6nZAM?vcYDg|+ey0NaYad4\\\\{-Ats/XVz"));
$write("%s",("b,roMmrb\\\\{azOz>aKl,NwJ\\\\}mtb<Gm1IdR=U:Ua7cd:vV45fs9\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'tnirpWMNga02(f\\\\{#LZQba4a4aja wohsn\\\\})8o3bo5Mqa904(f\\\\{#;)\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'\\\\})6307|5Tvg9439(f\\\\{#\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\',\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'&\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'(rt.\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'rupNaNq2:/r9P?|iWQagbTAFx7ev+1b./;+mbBE?aIyM<LOwCMsCaNa3zA\\\\}mQBa+exbwSybKA>y7F2/myI8ueybO\\\\{AaU07bJouqAagw=aBaCa=a@a\\\\}b@83r7c<+xbC:gbfR,bR42beb9bOaUax>LlW|S@wz\\\\}b,b0BY5Wp=I4bb=l<BaNyxo|uxT4b6beu|uxT:A5ntb<a=qZu,b\\\\{9scV3\\\\}wtbaGhv7s\\\\}pwz5B?arnMtW:f\\\\{|PZ62bNAU/R=|C?|-Bst=adthDdbYuN@5>s\\\\{Np8/J@jo5B?a/bS*6lp=8bm,Wa*b/J-\\\\}NAEa>a@8;fKyV.75OE2o.8abu5aIGO/nU-BaGo@T;x=.@wzvqnAJYaWa8vqnAJVU.oYn2<ZXdH4.1o.qabg\\\\{Cuym\\\\{FNa?ayb\\\\{pRWpPSns:=ayb*b/@,\\\\}4bSw6Bh|>yFwuI6b3bJ\\\\{s|k\\\\{0*tO\\\\}t.bG*+*<yY\\\\}rh>yjbjDlb+;o7.yat>a6SoA"));
$write("%s",("ttB|V/P:ko/b@avyVS7oVa?a;sAxi\\\\}AvXnZa\\\\{+13aRkhb/rr9YAwbl6tZZwnh,5\\\\{+rvZa<og@>a=axO2Qf5B-tbX1abd=k>VjxtEn\\\\}9*b*b6bc0>:EAPoM:ExYzvVg+OS-bs\\\\}@m<+qrtbB*G29s,x<TAa,\\\\{cmmsi0wwibabibq@V+Zq+bQ48bl-W=q.Cal\\\\{wUGt<?>/iA?7?@2r@0|OwnWad-|Z0pebXaZ:N@*oAa6.|b|0=25pQ9uC/*ab6?-w4N?XhZkZUaLpby\\\\},aItflbfboZGamZ748BVa>a5pZ:@3n<gJ7ekwI|iu,=,Ozb@T+;iHJyAa\\\\}o8;\\\\{SOa,qsz95wo4b\\\\{fjraz/-7b0m7yGp/bVSNa6c/**bM@ID@a|-I*ty6j+0R*R2K3NaZ.\\\\{tub<h/Xwb.@v+dbgbCrY5YjktzbEaDa|bf1sREGSw/lMl0yAagb*bCaP5qchbJ03bat,rl9vbFsW58boI6=LvIOjbA\\\\{y+q?7433dbZ7e3H-*u2n=0+Clb|Cs--bsJq@roCa.blb4bN+4bAa7exr5pp.UavcDa\\\\{+\\\\{b7bjbGu7,y+-wOaTlBaNa*bsJvbfByp\\\\{b\\\\{boC=;?aBvLTVdc>v0fbubs:4oP=UaL>O\\\\}ybm6H\\\\{jb7zWosJV+ub-b+bbb14;1Twx?7eA/\\\\}\\\\{+bX<O;|m>-ub3b:*2rZa1@VaJ+Ta+b-b,JnT+3VMEz2b+b7Vs@Vahb\\\\{\\"));
$write("%s",("\\}<av+fbVkGvtMtm5UYP>pb*7blUV/2n3bRa=yrp/*\\\\{\\\\}wmFaTVRVwC2b*bEVgJBaDfUFPa/vYu<2bbpNMmcR<a:-S=GTlb?a9P.bJo?d?GA/6b@aIyLmsy/CAVrlUaBwa8wb0/vL5z/n=tF7C|/LwbTa<ahwDTrt6UL9s?EScb\\\\}74Sf\\\\}RfQa*dMNxI|C6bZ0eb<m\\\\{,B+v/IxjzY?DokbAa93@=N5L-Eaz70uVniuLPVwUU3KIDVwYa1b9JSHG*\\\\}B8.w>qoP=53SaI5Q+GQc1(f\\\\{#alEF.fC?qUl2nH@;2ID5SQpop6oPqC|<0QpCaGannwG4>\\\\{3UaFxs-\\\\}biQ?.ebs-f<5-cb+Fr-8,e?c?gD*b7qhCebvbQ;@Db\\\\{ub\\\\}bZaSaItfbEr0yL+,bvup;|bG\\\\}Ya<tyb>CzoRzCuhb=KRaYuDTUaES*bAFFa,bCa7t\\\\{bN.rt<:7b?fEJZCizyFV\\\\}>utt+Td:/+mhiqePdqBm+s*IX=V=Sn*b3sT<aIYqGvSarpLcVdGa.CkbL.wbX=5b\\\\{bEx2,Gp*+lSgtpq-KRydS?vT<IHr9C0-t0b\\\\}7d\\\\{I4R37+wnv+\\\\}svKaw4ia\\\\{wo-bzbk<3bLoB|2n|3z3Jsw3MFSabLrJFI<2a</brxjbeb\\\\{Bzuxt6?mxO1|SmoOc-6F6TauSvKT-4bQ4Da1bGawD+bGaGxMu3z7e:txba5PaYaa5ibkboKmb5bi+/<FIFwrpLy"));
$write("%s",("myu5xp\"\"),\"& VbLf &\"(\"\";2ryZw=+*0fbrv0:dx4+0lFnLzMvrCYu|ud.==CwkbYat-\\\\{,tN9bP,qR\\\\{1TaRpgbgb/v9b+buvx\\\\}1b1b,be3wc>y9o-1w/u/uGXa-b\\\\{hkbs|R*>ay1/+V4ibGBgbEaWk4bQayb0PSorcv+rs+ea;8bJ0XojbHl2gBEZFPa+bXn7b/=lbAN?-tnc.<o*.aQU-/=Wb;Li3s;3bk.zQvcFahv+.k.=aTC,At;Qa<0B4w4PAmnp*wOfb0gY5?a\\\\},tn@a3bqH|.POy6vc@aYD/:*.1b>ISaN-vzR:D*y1@aP=?aNazC3L\\\\{f*bTa+2p*DuU-p|SEJ>ubU-.ukbCvU*4hrvVaWaC-f</+@FrEAL|rH*/b9qF54zVnAN9bE.*uub\\\\{p2n>:gbtbUa7bxbhzPqvb5>Z<rHYJi1Q:\\\\}8I8/bioF\\\\{gx\\\\{LnmR-tbovBE*blb*vdEiu2rJ.Catb6\\\\{ubgnoti\\\\}oqEazbsDxp3u+bT<Eobbbqkb*0Z01bm,U1Vtj,VaX@nqF8DaVa/bjh.Fyb65bsgbc.xO;.v\\\\}Va@FXamw=a|5Ral@F9I*Wa<o/*Aad9BN@NNa+/1n9>Znkn\\\\}xJ.Rf6y;m?J=|Nan9GCTM.bqnf/Rabb0=;+>aWa*.Ya\\\\}9LM.bPaUap2ul6b<=uyn9*o<4UaAao*B1a.Y5Ae,bhb5bGar/>3g<RaYnElTaebtmSn\\\\}bSa/,1t<a,y0."));
$write("%s",("@8\\\\{b=xwby,<2\\\\{b-ylnjz5bv+7bnr7bqhWl8DGC7ro8L:s5e@orbbS+DuvHdbxbsudE@aO1\\\\{b<aqnCtYwY5\\\\}\\\\{Ru\\\\}pFrh6cvIs-@OmOuQvEaf18tA1Y1so@aho-ds>Raj2kbxbZ0VxCaL\\\\}Lq>HWabbAaZDS\\\\{Va:c5lj\\\\{+\\\\{7babYa+bWL|K*v3bwJ\\\\}bF1/m7|Q,9pNaGC:I@<\\\\}bg*OygJM:atRyP5R-ebAaHJcm9E9b8B+\\\\{;2*oo+,yMm0+p\\\\{I9=ajbF0Ras--u+bNa,ATaV/<BHd.7p|6bEB<a,b=0hn+\\\\{\\\\{A\\\\{bVlgGCaTo7uH>Orlb/vhb\\\\}bd4R>H;6F9btsYa|b.>C\\\\{XaiqB0cEZuY5\\\\}b?aX2tndbWKqczb<aglhvXoVaGm.6GFPaPh65VrIngtj4YqSap3F0.p1boz,Kn3wbub<qVdum7F+\\\\{+ldbNoPqAF-bw9DaHJ6dp7.bmbjKD2zxeJzDl3p><ljxZaYr+>U/1bq,o,ubm,k,i,g,kb0uN?G9Qa9<tbS3O1J0o0OaFIJ.gl+I9b/mu6Pv6b*bw9Ua46L@S5p;XasqmtybyF\\\\{HGH.bRaSaCHs1.u/C6m\\\\{+kbjBv+Fa+/53n-d.nw\\\\{l9t=<ebBa-yg\\\\{9x-I/I-Ib5zbXo+IdHbb?p8zGa>?l,|bTCF<ibcb7b.bN5Ca/b>ICadrg*DIMIr6mbxy@nJp9=lb9/-d2tjx9/8pXwp2=I5"));
$write("%s",("BibVt\\\\}q\\\\{IyIb|2GD*fbBambYaRa0I9,wI\\\\{IY?Zw\\\\{\\\\}0t.I3oebzbab767bzbgl3bZwcblbwb,\\\\{5b.bgl@aGvNojxSalIIDE<GaXF0*FA<a>*c:i0lb\\\\{flbmb:ogtrCd\\\\{R-2b\\\\{b@,w>+0Ea1zhb8r./x02b?3v@,bLobbyw9sinZau8ybv+-y+doC7bNcUpPavb1EAa+zubub.6F-Uafs6?dbZs1h=aeb9<Va-bV.+Cg<?av:,yllkyFaKBmnUmCf>aNagu/@0BlbP8\\\\{lkG4pREtmiu5-,Fq6Zz:9leznF-e5bn3GCaq.\\\\}b-b/tPs-yf<a1v0Ho|zdbDatbwbcsxbRa2n.n3+Ba>0?79b|b3FJ+DxC7Baybl9bw.|EaEaLyzbmbDBFAIFwb,b+FprB0+l-b1>/bCa2w5p3p1b|-3bJ92xWaVawlCap.;+ab/n33u|m5@,5xw5?aWambk.Joeb=a0b7c9ranFohbAav+tbrl>y?a:4-oqANaO1GrElEaL+Pau,>a1bAwSa.b<q7qr9/b\\\\{/1bm3K\\\\}nBm/fw6bYEGn=lq+1lL\\\\{apYoWo/3zb9:j?2<m/3oZa\\\\}pp.Xafn75BzRahvGacqZ<tb6b?aH7,b>3yb0fwbPaD5>90fvw8bP,eb/qF88bk\\\\{=5Taib3uiyYACaYm6Azstb1lYB\\\\}b9<Hsf\\\\{fpztorY8J.6CRzZzXzW9B0f/S\\\\{;+-yTalbPDAafEabcpID"));
$write("%s",(">\\\\}MDS\\\\{kbzCM0KtlbEanCA6*oWaq::tw>\\\\}0/qEaGpFDv+Mu>CD@qt:D8DdxZaJ6/bNuT?UmJm7e|xGp8babCt4bXri30D,vg\\\\}mpvr1tybRq+bznMuvyKmGaPfKm7embdbJ1k.-b@oe,?+.b?l<amb8wybbb\\\\{b-b,bOa9bwblb6mgbVnabfbFa<2glysibV+Gtw0bb-\\\\}lbeCt;7qvbRa:-4-I?dt/v?a5bBaGaTv.sB|.bxbq@db\\\\{bL2ZvJsvrul-u7eCfTaR;Na-yxblb@s+bz;V2jbzx@aMl2wjbE.w;OazbZa53ErYast;2V/ib0;NBa/3moq9+-bI/2bvbNBMhq@ymF9upgbPaXaG/\\\\}bt;v+gb9<io2bWa\\\\{b6bq5y6:pT*twylcAWoPABag*Oabb8bzbhb<s<aN2fsRa-y+e+-vb?AzxHp9<,|;uG3RfVdY;VaF.Yz7y\\\\{b@aC0FA>aE.xqnq.b?.<2AoQmaq/bAac-gtdwEa0lLy-@462b,mPa|b74mb+eC84b75ibfbeb7o2pXkfb5bFa3nR\\\\{4blbZajr.bCaLr-@4/+:YuKl/@6?+\\\\{.bd\\\\{?,RfYl4bx>X2Dm>6Sz0=Ru*b/rdbhbjbtwqto;V>Yuvb1nPa@@1t5b>aS6Gp6bz>x>5h;=C\\\\{V/6b6b7e6c8blb.bAaTa7e<2v+BpE,tr2bImWlTaM<dx+:Ca6b+bx-Racwj?Dagbmswn\\\\{qxbdbbb4bTaGm33v"));
$write("%s",("xb5Z3C\\\\{e3X<x>338bL+rl5b\\\\{ywbR7ZrblPv8bTxp:2rtpebYa6o8rD38,BoWr/bF1A3vz7z,o1bW<rlcfW|Aa1bb|S60blb1w:-ubf2>0Faf?00/bOw-bovwbwn3u/bWp+>2br;0*\\\\{btbJmr;Rm?7ib/qzxI0Ga7.OaNuwn3bzbfq5vy1t/@=jby<bf<m?g-bUa1b2bSuC:Gaz<-okbdb.b9sqlazSkWaQ21bZzQmOml<1sMm3zibw4|bqm5:5ullIbAq?n,\\\\{0bPdFae50b,f3;BvEak\\\\{tbnqZa6bHpKz2b3\\\\{,d/bcb?ptb77Rapey<?aGaX+\\\\{bS;fpd;\\\\}bU=L.Zs@8muebp|tbfb.wllqnOa+bL-3oN+49SkBagbxb+bYaS2azNaen<adbEh-s-uubg11bub7vY7|nJ;Ju7rkb+b9=;m>aOa\\\\{bZ\\\\{abzbs1cbCa*bxbq2@albUaN<L<4b1bhz9tql0oO5xs=tP<\\\\}8l*!![2aba!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"g3b[2lpa\\\\})1(f\\\\{#(tnirP;)23&Z0/bgtJ;-bOaWoEwlqJ-A\\\\{=+Dau*SavzVaubk<zbP:7e;+-b/b=mRpOadfWa"));
$write("%s",("k|lb5z?vdbUar-7ek\\\\{G*2bhbSa0;l7v+,bEaxmr9abktibi04bRyb20ozv3;u3|b-<<+l,-5q+?fg<Nar;EuW:ebEaUa8pF:>0Ban<awabe*3/kbA:jbNaybvxNambVa*b>0scwbU/ps\\\\}bK;qppe2mdvdbzbUacw9bdbEopsBa5b6bvbEo\\\\}blbr;0fTaBy0oQa.wDa=akbRyGa-l+bCnAaNaXaMvs5cbfqM2=0>aPab-jbO7*be5fq-ykbp2e6lbXakbhb1bwbF\\\\{7/cb<a9sJgVl?fOq@0XaAq3yZa+b40B/7ehsCa3ba.3bhb?a2/mb2bcb24/vN5\\\\}pVa,b7b1z3b9blb3z\\\\{s+bdtQa1tl,Tarhgxjp7u+6Id1bZ.Wa4b4b\\\\}b,wgbErqpW3r+0bl/.w1bCa9+?++b2\\\\}P4zbHbguYq+bdb3p*b3uZ9vrIsAajbt5Pm/b5l48+blq,bdt,yOakbP4mbnrHxkbHlybwbyb/bTaF5:9Um8bGv=|dtPat.ybtw3bKs\\\\{2>*bbQ5fb1bLsr-+90n4b\\\\}pxtwbDo@aRa\\\\}bGnR*Oa\\\\}b3bO5J+ZyvbWa,qZdFa@vtb-o;+Om=2Yaf2otWaGaWmFaFvXasopf6bJ0Da*vwbs1+lR*K3F.EwOambebxeQazbtbSw\\\\}b1ldbmbF.DzBmGr\\\\{bmb\\\\}8fpDaz6m+zbrvxb1tot0+v+eqp,Z03bAaNp|m11-rf61p@a>aH3KhkyazYyVa7"));
$write("%s",("en-Fx*b0qG2xb9bVyY.l+QaPa*b\\\\{jub=ab1?v\\\\{2eb|pAakbjb+baqCt6bvpR*Gal1mb9z@6rn-b0/UlJ|QaGb:yqcM2fqB4*b7bz3fb83Mw8b\\\\{zC/e/6bYr\\\\{my6Qa*bKoirjb>aGzdbXaS\\\\{e,0g8bBa7i7bFaG+xmh,V\\\\}*0vb-rmb7y05qh-bPaab65d00z.ootf+dbTa3p3b\\\\{bV*csChDnhbY+5*tc6bRad/*bDaEa,b3b\\\\}b-r+rR*S/*0,pbb0oBrwb-.W,Ba7zHpjbFav+xbebgr.\\\\{?42bbbDa\\\\}b=atv,bSaCawb|bmeP,*28b|2;u0b2wDwGa@l\\\\{bRv2wCacbjbpq6b05Y+fb4byo5blb-bvb+04l7\\\\{\\\\{,zb=aGa@uflvb.rOvT*6\\\\{Ra.b=aN\\\\}Aw/thb?2jbdbD2WaQaDs0zAa=azbSamb6tfbWa-u>a**|*@,1bk4gb1\\\\{Ta,y3b|r8/?aBantQamewlFae3Uabbhra,jb7bl,\\\\{/5bhbL-Va9p*bbbgb0b,bqooo*tKt0m6b*+D|Pa6tNc4.bbF1vchbFpabSaebhb<qFa/b||Waot@\\\\}XaVaFxabMqGr|4WlqtFwk\\\\{bs>a\\\\}l-+7e7ecb0bqnv+iba/7eMql,T-mbcb5*yu1sPaC\\\\{cbX,8rcbybQm1x6\\\\{Pa;ykh2,6nQ1Aazbvb\\\\}\\\\{cbxbNx.b1x4bvyxbDa,d\\\\}b0btbO+kboza.7b"));
$write("%s",("8bPa5b>hf\\\\{Oap.?avyOompVawoyb<tPaDp5nen?aQay2ubn3R2ZaHqlt*tApm35ncb+bWr7+frib+/;0\\\\}p0bDaC0+bN2Mp2b>a?s.bAoEr1bkb=nopZ1kbfbzbtsfb=aT*\\\\{b0b|bmb5*3b,l-mZaab|b/bUaYarttbcsqyvb0b/bpqbsXlJt7e\\\\{bRatb6,1tWb5bib\\\\{b|bpr6bZaK/-.UaxbZa1ncbgb=irzybNaK|:pTav+cbPtwbRh/bDpQa>aHq-bybVnmbOavbjbubVl,yo\\\\}xbPmt-ZtTaM\\\\}P-8t,b=,Z\\\\}Vaapt|9bTai1xs+bFaP/0uJm5zKoDa5b4bm0Ta5b2|Fv=+abgbmbPaSajbRzGpUaFaRv9nYav/X*7eTa9b<y0b8rbbtbI*kbTa8bvbgb,b6\\\\{Zo/beb0fAoGqsqg\\\\{Xafr4bh0kb3bjb30jb5bi\\\\{kb5bZaaf0b//OaxbjbpfWofbYa7y?xhbub8bxbs/jbmb|+Wx0bbbmb3b0bu|Qa=aXa\\\\{b=a9bcbMwwskbgyl-rvSrgr0b4bPae*Mq,mExybdb2,1w7bh-hzz-wbNa5lab0fxbtbBav+ubtvxb:t=a4bbbabjmtbYavbzbhzu\\\\{0b5bTa1qSa=aibhs-bNa@afbfbA\\\\}PaZa5bCt\\\\}qzbp.tx0.OaupcbJoDa,b=amb7e.bh/:z6wdxubabRmS\\\\{?fE\\\\{EaTaub+,=xJtcb*bubxs7b3b?aYa7"));
$write("%s",("b?nGsUo*tbbHq6bPa0bxb+pWdcbzb0*ab.lFmUpeb6v4bqlWajtov7e5bUa2bPaCa\\\\},;zubE,7bkbWatfVaj.|bEa,mm+=w5pUa2gRa9+vbybRa/|o\\\\}Xawz8bSaU-+e:-tneqPaVa@aVab+7eWa8b=-gb?a3uPa+yVpRx3b7c>aEnwbvb>amxhbTaSaVambtyc+suDxlbVq,tPaWav+0bublb3baq?uPafbRaCrVp2t5bQacbSa0bFaPa>a-dg-7,?aPaibDn?|7zDaebtblz:lin/gab1nYrCa,b<av,O\\\\{Tm\\\\{b7eP*Om\\\\}n3o+oUa.b7,\\\\{z\\\\{fHoi*GqH\\\\{P+\\\\}w6*xbJzi*?,dxjbQa/vFal\\\\}fbcb.btbXaAaRm.,.bOa+z\\\\{nOaablc;zEw>l3b9tDadv>aTavbVa9b9tey?a<a2bvpOzBacbmh+b2c3blqMvwb-vncAa\\\\}buc7ewbY*8b|bKofbswg\\\\}=a\\\\{bebhoib?vtbib+h\\\\{fWq/bRakblbzb,|fb|blb2bDa8bAax\\\\}\\\\{bDa6dZabbTa*+jbabvc>aSaxbEaBaUaEa,wfbhb4aU|Ra,bYkjb4brlEatcgb<ac+=avbTw4b5bjbJo3b@atuNa=a/b\\\\}*SalbkbEa4b,*;x\\\\}*@\\\\{z*dtSaTaWaAaSaAa*uUaTa=aZwG\\\\}\\\\{bgbPx+zRaTavz?a0bTaUaHd/bkoGdVaRa2bjbglmbmwEaab|r@a3ugll*"));
$write("%s",("Wa=anewtuytywzSa@amb@a\\\\{eQaXaGaiw5p,bBazb:\\\\{+b9bBamrDf\\\\}bubNxtb7zqo4bXatbeb,b2\\\\}Lymbq|hbNpwbSa;q9q,bbbswXa*bzzCa?aib,to\\\\}FaYa>qRxtbXvWb3bLrbb/bNlssZzFv5b1bYa6bPteb8bUo3b7zjbSa\\\\}bZpDaWa>a8okb3udb,b9br|:p0oFaZnKt.bFaXh=z+b:pM\\\\{K\\\\{I\\\\{e|F\\\\{D\\\\{Aq3pRa\\\\{bb|unAaeb5bNa0bGp6nlbeb\\\\{b0wCrmwBp/wbbdbu|Yrlq3qxoF\\\\{DaRa.u-b9b<aPqtbawRvlbtbnr3ytbVrmbabOmVaXaF\\\\{Mukq3btvOutbVaH\\\\{TaUnZzXaAt>a8bPsFaRaZaE\\\\{jb<auq9b\\\\}b.o0z=aVajb=aCa0ltbaboqkb2gabWa<u.\\\\{VsioWadb6bzbWaBa@acr9b;m2b8bZa9bp\\\\{Qa+b@a,b6br\\\\{6mwbXrVr\\\\}w.bvbNawb3rXa0bvbZtEaFadb>a,bFa?a/qkb:z@a\\\\{bwbWaYqNa7b4bfb\\\\{bAa7rub7b7rRawb5bRw1q*pXa.bkb6bZuzb?x=n\\\\{ugkfxtcmb1b=tab4bUacbswxbxbTa-bkbqq+b7yibNaFnAa5b5bzbooVaTaqwlbRa/b9byo7bjucbubTabbcbbb<aYa?aDalbhbkbvbhbHr@twb\\\\{uop/bZa-y+y3y9bjbUajbybDaBaeq.s.d2"));
$write("%s",("bYn4b7bybrs|bTaZa2bFa0y0bZaUa,y*yfb2brh7e9oUaNa8b\\\\{bjb;mDaVp2bJcSaPamblbVaVaOaWahbcbQpEabbubyohbJgXaFr2bcw8qUagbtrVa|b6bXaTagbjtWa|b@anr=aabRtPtOm\\\\}b7eYad!![2aba!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"g3b[2lpa\\\\})1(f\\\\{#(tnirP;)23&=,b8bEaJcPt3bRqOa*bPaQq.bNuRambGanpSaXaRa8bib:cFmgb>a5b/bRv2bSaSn7b/b3tDa3bDwtbOswb3bErqfGa\\\\}czbzmubQa4ack6u|bWaRaVaAa@aSa?a\\\\{bWaNa,bdbEa8vbf7e.vtbAeybNt5bSa,b*b/btbCa4b*bNpkrbbWasoYu\\\\}b2bZaBa.bwvFrrqmb/b0bwb/b=aubzb-r?a2c:v8v2bgwvbPaWribEaCaWa\\\\}b*b.bVa2bGl7e3bZacbNaaptbmb|bNa-b\\\\{qdb,lEtmo4b=seb.bibtbkb7b*b2vBrdb6cXacbJgctQa\\\\{bTaTaQaxb?acbvmCaQa8b6bkbkb@d0b\\\\{vjm0bPaToabTa6dbbPlNp2b7bwtjhwujtYafbjhCaCoWaXa"));
$write("%s",("mrarBa3bwbvcEafp7ezb/bBafbWkkbQaWkQsmnqoPaPa\\\\{b.bUkYaab0bWa3oQaJmcb\\\\{bib1bQa6b<a7eab3bBa>a.b8b,rZa4akpPrAa3buborwbUa7o@aUa0oOa.b.b4bRa1bktSqQawbcbRaRatlGqaf>aqq<aSacuWaUa8b7b7bVa4bhbeb6o3b7brt3babirbb+babmbEa;q6btb:cibzb?anl-b>h7bYa9bXalbEr8t7n@aDaFrXaXambybgb7bnofb8b+bBa\\\\}b\\\\{b2b1bTajbxbEqYajb4lTaBaOmFsybcbOaXaLrEafbbbZamb=aWoCr.bdbooYagb|b\\\\{b1b9bRa9b0b<afb3c\\\\}bkb/bwbgbmnYaNa\\\\{blbvbXagbZd\\\\{bXa|b,bNavb<aCaFa8bHoZa*bcbBa7o\\\\{bksbs/bZl+b,b;m5hFafblbdbebjbAaBaebmhbbbbNaEa6bNa?d|b*byb7e6bKlYa+r+b4b;qFaOaFd|bRaubcbEa*lxo\\\\}bPaqmip6b/babXa9phb@azblb7bvbDnwb-b>qibNpJl4p,buqMpAatbdbkehbznub7eRkRlgb\\\\}bwbababcbWaTaybflwb0bDhYaRn7eEadb-bmbBaabvb2babybQa|bCadbYllb|bOaubibgbZagb4bZaVl0f\\\\}bmbZaubkbmb0b6bxbylbbzb7bOadb:cWpeboleb\\\\}bEatbgbubAa>afbwbpqdnYa3oBa/b2"));
$write("%s",("b\\\\}btb7btbfcSaVn|bKpep0b-bgq0bEa0b8b/bXaZa,bUocb?aZaFaSaOa|bkb7e9bvb,bRa?pVakbgbXa:c,bebWa6oKpdb|b7b0bRafcXaabxb>hVavbdbYaTkNa.bboJc\\\\}b7bEa-b7eVlY\"\"),\"& VbLf &\"(\"\"abbeb7eRa|byb@asm\\\\}bzbTaFa7bSakbFa>aJmFa\\\\}b@all5bwbCa7eibwbXhVhekqm*bKnZaWaJl?a\\\\}bdb/bSaubvbeb0bkbVa5bLh<aTa|b1nibTaYa.b-b\\\\{bYakb9b.b?aebFazbebQaSa\\\\{brcVaFa*bzb;mabQaUa/bvb7bmbmbXafbib0b0b7eybXaUaOaEl5nQa,bTaNa5b3b,b7eSaQaYaFa|b|ndoyb9bPaybTa1bFa.bXlebSaVmfbEa8bgl.bwb*b0b7b\\\\{n\\\\{bPajbwbkb8bQaub0byb2bafPaHbvntnSa1btbjbcb9bzbjbRazb2bVa.bXkUa>lwbRa0bab\\\\}b1bdbcb1bUaab>aQaZmXm*b2b|bUavb@aYaEavb*b5b*hZa7bPlwbQfQa1b-bab5bDaubtb|bDaUaPa7bDa@aFa1bWarl6b|b<aFa+bWa,bzbOa,b5bcljb|lhb*bBaDavb+hcbmbhbvblb7e>a*bjbhblbYaZa-bib2bXavb4aomdkfk2b6bcbRh>ajbDa4bNaDakb=a>aKh*bAaFambwbzbdbGbjbPa,bAaYayb4bub>ag"));
$write("%s",("b@a5b,bvb6bab*b7e7b<a>adbfbefYa5l|b4bxbybPaGijbTaabFa7e1bebibjbjb-b5b+hebPa7erl-bTa>aFalb,b0b=a7bdbCaEaybVdQa4bSa>aDa*bibBadb9b*b-bEa7b6bAaEaKk.kSi6ipkkkAkGi-a+jNj5kZhai/k9kFdQilk1k;afiykskRioj.jYiwk6iuk\\\\}kzjLjxkdjCaCeMjjkwbXbNi>jRjliji@jSj8jEajitj-iHiFi3j?jKj@i4aWhbk9aXhHfUh/b-b4bCeEfub+eNi+jEj7jbjdhAj-jZd=jhi9aEa.i9jxj0j-ahg4jDi,juh*jwd:azjlj1j=aAaojuj3iyjejkiajPimjPaxhkj<g<a-bfiMirjjjaj5iOifj9i+ibjMfZiNidhLicj:aCaaiCiTi>aAa-a*f|iIi+i9aai:i,iAaEdxfEigi2ihgBizbmizi8iBaCe4iuiIh0i*bNcsf-d5bxbfi1inixi@axfii\\\\{b\\\\{ipi*fsiOaaitiyi?aAaxfviaieimiFajihifioidi9afiHaSeSh8aCa@aCe1b+d8aZhMe8arb8a8a2b4a4a3aGf4a-exb3bHb6bxfCgzbxbubHaMfFgreIg3b4b.b-e,cCe\\\\{c1bzb.b1b\\\\{h/hvhthNg?a=aGf8btbhhthKfRgzg>aBamgYf?atg+gOb\\\\}gZdobfhogBa?amg|b|bvbaf.b3b>bTdObchTe*g\\\\{gcgEdmgzbIb"));
$write("%s",("Efrb3bzejgegrgMfpg@aCamg2b3btf:b*f7fSeQeIb:cCewd-b3a?a@a3aKa\\\\{b;apcwbxeIa3b1b?f,b|b0aTdZcWeSbgghgsgHf@aagBe@eTdYcJffg*fdgBaGf-eybYfXeNf5fLfreSeIfDa3a3fifOe1aEc1aSbRbubwb7e,btePa/eUe*fRe3a>a3a1bxewb+bxfPefc/b8b1bJbxb;a:bSesdZdEc.eSe<e;cZaxfrffc5baeVewfoctbxe-aSeNd6c4c/bCewbAe3b|c;a<bre:bre3bCe8b5c,bxb2b2btb;a?aie:eZc8ePa9e3e-eJbvdHareKe6dGa6exb-b6c4a-are.b\\\\{bmcMajare-breZddd2eGa+b-dtereGa5aZdYc?cre4c2bzb;azb-bHb3b2bJa7b?aSdaeYdRaYaOaVafbVaibTdddRdPd-a?a;a>a-aPaBaedVaNaUa?a?aed-aebcbkdvbpbEabc7b=aEaAa?a>anb-dub.b+bzb>bMa/a?c9ajc<bFaFa9a>a:b;ajcIc+b+btb\\\\{bvb3b:c>bYbWbjcKbIbGb;akd6a6ajcfdedXcadDcddCbbd6a/aZcddZcCcWcCcYcEcjc9a2b5aOcMcKcIcxbvbtb+b/bxb1b5a1a/aEcSb/aObic9aCbNb:aIaIbtb,b:avb|b+bub4bcb-bpcnclcHaebdbJaGaxb,btb-b8a1bxbwbtbxbUa-b.b|b3bvbxbfb/aSbnb5"));
$write("%s",("aIb.b\\\\}b-aIb-avb-a1b.bybHa6aCbObsb*bCbobBbNaHa3b-b|b1b/bJaNa/aob5a/a5aJa2bg[~ia3(f\\\\{#,43.3\\\\}ia9541(f\\\\{#X3~ma(f\\\\{#(tnirP;)23\\\\}ja7362(f\\\\{# [4Lma5904(f\\\\{#q\\\\})6j3bh4Tg5Mda132g7Tja5683(f\\\\{#&[2iha=s,y=z,s6[\\\\{8Qea0603+:Vba0-;\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'i6[Y3+|8jk5[-;Hba76?Uca560<a7>[u8[6=iyay,]99999[gnirtS wen=][c n3aea\\\\{)v]y3b&a(niam diov citats cilbup\\\\{RQ ssalc[4Lba7@DVea9493$?[h9Uba3~@Wba3~@bj:[9a& cdln&&&&;maertStnirP/oi/avajL tuo/metsyS/gnal/avaja:b&ategn&&&&2 kcats timil.n&&&&]; V);=:a;3ecaL[I:aD:hha dohtem;3a/4nga repus~3acaRQ83cgassalc.|>[\\\\{:Rba5>E(\\\\}9-ca14#:(i6[\\\\{:.oa(=:s;0=:c=:i;)o9ajaerudecorp>=Mba0$Ma>=Qba9-R[PF[g5Qca75.RUza1251(f\\\\{#&(tnirp.biL.oken\\\\{,9bianoitcnuf/G[96[A8[.3cba1BNWK;[qa(rtStup=niam\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'tni[>Nx8dkawohsn\\\\})840h;\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\'MJ+ba8~7Uda332Z4Qea1918c@Xha=q\\\\})486h6Uca148GQba7f9bta(amirpmi oicDAx\\\\})42QIaca3Cl3fpani;RQ omtirogla?9Ml4bk6aea.tmf>Acfacnuf;t4Tdatmf[3Ugaropmi;|Jafagakcay>Mda115)6dbapu6Mc4bba-X3Sjatnirp tesu=MyIaca(n)BQca725:a#a,s(llAetirW;)(resUtxeTtuptuO=:$5Mca36)6ea4RdaS CZ3M.3aca&(X4Rba [5[[5SiaRQ margof5O.3ajaS D : ; Rm5Tba\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'X3Sqa. EPYT B C : ; Aj5Tka)*,*(ETIRWt5UhaA B : ;e4Sba [2cj5Vba:a4(+3[+3wda(nfKC&;Ya|a(etirwf:oin\\\\})8(f\\\\{#>-)_(niamp3cpD~ka(f\\\\{# cnirpP@~T4ahastup.OIVO,FLataM diov\\\\{noitacilppA:$[cea[06xE3k75a*Mcpadiov;oidts.dts 5Ka14\\\\{kaenil-etirw45lva(,\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'s%\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'(gol.elosnoc;)\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'K3s[2cya\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\' nioj.)1+n(yarrA>-)n(=ff4kia!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\}54,1\\\\{.n3cja# qes-er(YRdba&l5rba!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"$Sk$3lo3r33tla1% ecalper.S4l(3cs=gsarts(# pam(]YALPSIDq6cua!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\".NOISIVID ERUDECORPU3kma.RQ .DI-MARG~3oE3dnaNOITACIFITNEDG9dsa[tac-yzal(s[qesod(n6apa!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\");\\\\}\\\\}!\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\");\\\\}/****/e3a\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"),s[99999],*q=s;int main()\\\\{int n,m;for(;*p;)\\\\{n=(*p-5)%92+(p[1]-5)%92*87;p+=2;if(n>3999)for(m=(*p++-5)%92+6;m--;q++)*q=q[4000-n];else for(;n--;)*q++=*p++;\\\\}puts(s);return 0;\\\\}\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\");gsub(/!/,\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\",s);for(print\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"define void f(n)\\\\{\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"00g,\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";for(m=1;m<256;m*=2)\\\\{\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\""));
$write("%s",("\\\\\\\\\\\"\"00g,4,:\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";if(n/m%2)\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"4+\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\",\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";\\\\};\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"4,:,\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\}\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"389**6+44*6+00p45*,\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\"));
$write("%s",("\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";++j<=length(s);print\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"f(\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"n\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\");\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\")for(n=9;substr(s,j,1)!=sprintf(\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"%c\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\",++n););s=\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"4,:,\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";split(\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"145 160 17 17 17 23 252 141 0 46 125 231 229 231 250 151 243 243 243 231 231 207 159 63 4 231 249 255 191 225 17 127 206 103 51 57 152 37 255 57 204 230 103 48 79 159 159 151 252 231 51 51 57 193 47 249 204 230 102 115 4 251 190 249 243 207 57 206 115 158 9 231 57 156 206 102 9 193 48 96 22 236\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\",a);for(i in a)\\\\{s=s 0;for(c=a[i]+0;c;c--)s=s\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"1+\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";s=s\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\",\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";\\\\}print s\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"@\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\nquit\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\"));
$write("%s",("\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\}\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\")');\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";FORiTO UPBtDO INTn:=ABSt[i];print(REPR(50+n%64)+c+REPR(50+n%8MOD8)+c+REPR(50+nMOD8)+b+\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"J\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"+a)OD\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\"\");end;\\\"\")\\nsys.exit 0}\"\")]]></xsl:template></xsl:stylesheet>\":s=\"   \":For i=0To 7:s &=Chr(32-(Asc(c)>>7-i And 1)*23):Next:System.Console.Write(s &n &Chr(9)&n &\"  \"):Next:System.Console.Write(n &n &n):End Sub:End Module"));
end endmodule