module QR;initial begin $write("%s",("Module QR:Sub Main():Dim s,n,i,c As Object:n=Chr(10):For Each c in\"<?xml version='1.0'?><?xml-stylesheet type='text/xsl'href='QR.xslt'?><xsl:stylesheet version='1.0' xmlns:xsl='http://www.w3.org/1999/XSL/Transform'><xsl:output method='text'/><xsl:template match='/'><![CDATA[write,format=\"\"%s%s%s\"\",\"& VbLf &\"(\"\"\\\\write{-}{txt}{(\\\"\"with Ada.Text_Io;procedure qr is begin Ada.Text_Io.Put_Line(\\\\\\\\\\\"\"print\\\\\\\\\\\"\"\\\\\\\\\\\"\"STRINGz:=REPR226+REPR153,a:=z+REPR166,b:=a+\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"2\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"+z+REPR160,c:=b+\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"8\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"+z+REPR165,t:=\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"write('implement main()=print(\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"BEGIN\\\\{s=(\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"#include<stdio.h>\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\nchar*p=(\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"Ra#include<iostream>!nint main()\\\\{std::cout<<(!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"class Program\\\\{public static void M83apbSystem.Console.Write(!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"let f(c :Int):Latin1=if c=127then!!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"!!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"else(string_of c@!!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\" g caffeine !!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"@$3kEa!!!!n!!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\")@f(c+1)in print(!!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"Quine Relay Coffee.!!!!n!!!!nIngredientsq3aha!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"@f 10U3cgaMethodz3c#a);let g(String ->[])!!!!n[c;t]->w4edaPutY4spa(int_of_char c)05auainto the mixing bowl|4ejag t!!!!n|_ k4gtaLiquify contents ofE3oeaPour\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'3w\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'4elabaking dishv6biaServes 164doain g(!!!!!!!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\")))s!![2aca!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\" [2bo3cparts(nltnirp(])]v3cja.NUR POTSp3cx3dp3jba!!M3dp3df4fda[))j3ci3e,3cp3l[2kga\\\\};)06xu3kgaqp]\\\\}\\\\};@3\\\\}ga)1(f\\\\{#+3~ba3+3&ga7(f\\\\{#.,3~ba5&4\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'ga13(f\\\\{#+3O97l,3tkaD ; EYB RC73(da,43.3\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'daDNEZ3Sda. Ab5VeaPOTSc5Wb5TmaRQ margorp dS@aj4ObaSj5UV3Lca36V3Vba&P5MX3agaS POOLi;Vea\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'&,)i;Uga. TNUOf5Tfa(rahco7Nh5cgaB OD 0l;Uca&,t9Rca)At:Vo:UiaEUNITNOC0Kaca01l4Mba7\\\\{>&ka(f\\\\{#(tnirPJJ#ca52q9aj9Vm8OxCceaRC .b4Ska,1=I 01 OD3GWcaPUc4Tw<Rva;TIUQ;)s(maertSesolC;4Rm|;=ka21(f\\\\{#n\\\\})8i3a"));
$write("%s",("g4Mba5*;aX3Mia115(f\\\\{#\\\\}Y3Mla3201(f\\\\{#mifEU$g7*da402h7cj3bh7Mpa904(f\\\\{#;)\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'\\\\})6992:\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'A@-da983w9aka\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\',\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'&\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'(rt.\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'(7Oba8v6\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'k5-ba30;b=>My7ceaq\\\\})6j3bh4Tg5Oca51h7Tca101>aca\\\\}\\\\}2<Nb6Wj8[ea\\\\})55#=Uea1473h6Yea&dnek8[w?Ica02c7Uda398l9[t;[$a\\\\{#&&&PUEVIGESAELPn&&&&1,TUODAERs3a$4Lda938<?Uea7522:>[-8[g5Oda116@WUca84BVa$a&&(etirw;\\\\};u=:c;))652%%)u-c((||\\\\}6[)8Qca00+5a5:Qba9.7\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'h6[T>.da#-<b5[CSGca01\\\\}PUea98917>[l8[ia\\\\{#&&&||iz=Nda158=?Uba4vIaEC[m8Qca76$Nax:Qh6[la&&&#BUS1,ODv;[p8Sba4/>Uda106iL\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'i6[q8.WHbma)3/4%%i(&&&&HT[Y3Hca31zPUea16924>[\\\\{OVba5W4(=B/\\\\}9b/UR\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\';[m8Yda197/?Uea50311>[.TdNa2=:/t;2%%t+2*u=:u\\\\{"));
$write("%s",("od7 ot0 yreve;i-=:u;1=:+i\\\\{od))1(evom(dro=:t elihw?s;)s*iU[iUTca22$?Uda778i9\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'i6[jU1HIQ\\\\}@Wba1p9[(D[vXQba2k:(XP.ba6o<aHJfi6[q8[h4Jda955$?Vda352&>[nb&n&&&&dohtem dne.n&&&&nrutern&&&&V);gnirtS/gnal/avajL(nltnirp/maertStnirP/oi/avaj lautrivekovnin&&&&u9[Y3Fca32*@Vca37u:[\\\\}<[da\\\\{#&[2aeb\\\\}\\\\}\\\\}\\\\};0=q;)]q[c=z(tnirp.tuo.metsyS;)0(tArahc.y+z=]++n[c;y:]q[c?n<q=y\\\\{)0>2%%++i(fi;48%%)31-)i:3c&as(+87*q=q\\\\{);07951<i;(rof;n)rahc(+=8Mca42bBUda358xOZ>9[g5Rca10>ZVda803@:f[2cm6[u8Qea2783>VU&;(h6[U?2[2coa=]n[c);621<n++L>aqa0=q,0=n,0=i tni;35[CJGca93S?Uea7961T>[=8[=8lfd6a2b9a4a2b2a4a5azb@d;axb<H2bqcvbGa6aUcYfLa4aqc0c-bat4aJaJaYf-ayb.bJq?*Hagdgdrf;fHawb;f6apb7b?lnbCbTf|bUs;dLb>aSi2a6a|bKaKa6a2m:a@aEa2avb5a5aveHaAa\\\\{GV*JabcXbVbjc+hDh1BCf3bo|.dE-JaMa\\\\}b"));
$write("%s",("JaPaCfwsJaJarcJaJaTaJa8b+B;a8bMYKao?k|ZKr\\\\}vRSaQ6BPKa8bQ6?aTao?o?k|Nao|\\\\}bJaLaJa8b@*Nah4cqa8bNa|U1B:b+b3b+b)BQea(f\\\\{#\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'5agar\\\\}JaHa|4a<4a+aHaJaJaQays;a8b1O:aUa:a+BCb2fbcZbXbVbwbk7gea>a8ao7bnacohlEjc7aCbTfu7aoa+i2a6a\\\\}bKaKavbg7aXa=aMO:aGaCaJadczdUbCcohjc7aEaqbCcKgsbsb;dLbTb2fObldidpbjcHagdidpbrdCc8d=a-a<gbc3bJcrm3bea|b9ai3fEad7apbX4JdHdRihcye/bJb|cs\\\\}RhTV7aX45a2bIgMa<gbc.d62Ja>a2a:b6a5a-bBy3biaGeU/vc6a53kxbxbA@i8vckd=a=addqelbOa-aRalbOawP7RteQdfeteGh7b3f|hMiHh*f.f;fGhEgKg-ewcef4b-bjh9a4aSeqgig7hTh/bJc;a\\\\{eWgCe\\\\{<NIJc33aO;c/a9aWhGh|k2a-eepGhte>jwh4aMiHhdh4f*fZf6l0bMe\\\\{3c*bMf-h8d*fZfJcGhXgyeUcOkQhjbC4\\\\}c<H=v6U;a,bRhHNfbpbreub6cXbvb|@nbreCeo0,fCe.d62zh-heh7hVhEaEdajAf?g=gHf9a7btcCeyD\\\\{l=g3a=a9a:Pxbq3e33gea3aAa53icaHf33kha,b9a7bmW3f%av"));
$write("%s",("yBa+h9a7bUWCeyD,b7e2g+-Vg-b=g3ak3a1aCe+bBd@d\\\\{e=g3asb>gAa3aMeGhXeqgQghgOgbg>gEa3as3gcang.6coaSeqg,h;glfMe=a-7cE3icaMgA3bqBMxa52(f\\\\{#(ntnirpn\\\\})821(f\\\\{#~>#n40\\\\{5blbs=GfGhlf7eGgZfdp2b2a2a9uThkg1i.f;fMeGh-,8aGhpbhgHh*f2fJaJaubve3fKgCe=anbre3flgyb6g-e,bJaGh7b5a*fZfI3cA3esa9a9b9aMg3flgCeGh>aq3acatuq3c-a-,:a|b9a0b9a-,7aGh-,Ia|b-e:a9bJa0b3flgBjS3c%aMg9aCaAaJa9b3flgnbreJaEgoh-e,bMem5g1a3fKgw2CeDdMfidpbrenmCenmCeEggf-eA@+dCenm.Jbbw3aeaGh7bw3iqanmnb*fDg\\\\{f+sJc6a24a0a8b9a7b-eMaJayb>aX5cXJa|bCezdMelfjfJa\\\\{pcXJa-s3b,aGhGhrK2b-e+b|bOc:a+hJaub-e.dOcbm4b-bJa3p>jiashqh3a3b.>iZ:aoa*h3a.\\\\{Ge=g*h3aT:e6j5h3h;awb;fGhnm8+-d<iHaJkvkEkciIi-k+kEkNk/jLk=k.b;rMq=aI@Q?|.N?Nx,b7e=6,bGa7J2g39v01sA?QY1CXGCazTz23xY1@GK*3xzbjtF*;tMpM:HIQtb3x*NlH/=acl=lZl=aFaN,k?XGNlgbTp2b</Ta0zU=>"));
$write("%s",("aYa<;Daqrx*lThrkbX?*yvbcb@a8Khb\\\\{nAa\\\\}GEaC:nsD3k7Ba-9;y0n@|T7WaKmmb.ozDl|lbSa\\\\{XsvEaCaDak?cyT+/y.bHL,/DZgb8Edbrr+mqq1R<yPam/ItlF2oBxlbty;3cnzpyya7-bS=\\\\}t\\\\}pxnyFHqh1irD.Gr\\\\}p?\\\\{nK\\\\}N|+v7s8NrhbBnslonT@ZQ?u3mAV/,YGib\\\\{XMquwNaBKp\\\\{Yx1blUDa?Hq.hGSa\\\\}rab<zB0n4no/b\\\\}N;0/bWaFaItSs<h+mF*Co7\\\\{ZK<H\\\\}IEn\\\\}7?m,b0z\\\\{ngSR\\\\{M1R+J53bBxtL/tmbAv=/Z/6VJTbbwbq*g64*VoCLh|>a\\\\{7h<OGY\\\\{Da0t8bXaA0yK>zOa@mkhvbhn@J:cR\\\\{ab43W@Y?ZSdbyb>aLSIwL|Mq8+,bdbu*|vvbF1Em@n1n0fSqIJ2bXsT*7*B0ly;RyDY|DwLvUs/b8tdbEoHI,b?nVdmL,bf9<abbq-dlx.3v<4YxKlo=iA2@Klhb8mj\\\\{Fujb2bE=3blbDau9k@hb6b+r==KlNaYarLhOeRyGLr1=SarlO9,=*=|=z=n@Waw=7*DarrBNzbg;=Ds=2bw<?pqraOpulbOm|PO@noaOZ-Da7*Dah,f,=aOaZrBaXaCm?;j+37wzwlkbMYpln3Ya/\\\\}jbJ+n3oB=a?ae3au3aaedMOaUa/<Sa,b1bUFtN:\\\\{Gs1<BaEagbCynK|<A=6b:Jw<,b"));
$write("%s",("2</mZaPs:JpxUKE+dlzphRY:DGdblbg<=aa<jl6mBaEa5s0|lbkZnrr+VN7yQ,vCDNRzEa\\\\{bklv9\\\\{RYuSaEo|by+EaH,jl0m+y8;nrzb;CK*nrNaav66i\\\\}cHx*lEx*aYBafb-wmbDa6wjl0/aO\\\\}WEa0/Pq-wWaq;qUoBMvYa/\\\\}F4pvyyQxk?2bH+Rn,->=W9AN\\\\{8DaNE5mMML*-=auP:ERTabN.mzo0bCaoFR\\\\{DaPAYkhbOnDa-b>36brtpt7bgwk0\\\\{nllhbl*qs?\\\\{23=l;l?aDPV\\\\{+Bhb<ADaR47e.8KrBKs=m3a\\\\{aDa-b2mn:l:hb5hDa-b:;f:Mxo*%3cvbT*MxZl@aOaDa@\\\\{nqhbu<qZ\\\\}Hmq=a+Bhb<aGPKLq:ebKon>=@z*Yau\\\\{D3Da*m*bDaW.6bYsDaR77b3m|bv9bo@p=a@7D3+m0pBOa.g<4Uz2tm/3icbF=,5d8jbPCCYzADa:cDaPaEG\\\\}I?FRBg@KBCr<a2m=@sFebq?4w>aKmYlKplb;rSaF30bYrxn?x2mOaeV+yhb548+Nk3b=dbF-9=l-U9qMqmb.wHz@aym<arImFu|F30baPAaY.Na4b\\\\{eqDrrSqvoZa62zpD4mb,b<|kqWNCa2b;;20/bYj54M1hRhuXvQXvbn@I4qltqBa4bJ@H\\\\}>XvlTo4b;8@I5z+b?pFrzmto>ahMub\\\\}byKhN3b5qcy**f4VaDagbfn2:z=Za7pxbu\\\\{t<"));
$write("%s",("KqmbBxbbOmhbub3RnlLcCxxbwCeUH?;9cNL7It0bJUWxjU>a*b@u+o<u1bDaY1ub?/\\\\{f>0J4Fa<aw29.0;=a+yqUC9e2G+>pWaBwOB\\\\}bNa8+|vqtjbWngGGa7JWLgb+/K\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'tnirpWMNga02(f\\\\{#LZQba4a4aja wohsn\\\\})8o3bo5Mqa904(f\\\\{#;)\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'\\\\})6307|5TKg9439(f\\\\{#\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\',\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'&\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'(rt.\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'\\\\{@l=rb2t?OwX8zD,r<HQ\\\\}UsOt\\\\}6mb,bfAlyI8Mpyb8.Eae2Nae;\\\\}<2?7bX8=a@\\\\{|m9bi9;yAaw3QuCa>aQWQuvpGaL+2Mt9VasU34:vXkWk@32MVMLLhQ\\\\}zFaSA.8yrxRr=ypqteuk\\\\{|bxzdMU1zb3/g.7n2v?s,b5bz\\\\{Wb4balUa6FWsYaMq5bcFh7XGCaTI,Q=.zb7eYpN\\\\}\\\\}n2bg.,\\\\}kboQT:fVNajs=a3bor\\\\{*QwfDamz\\\\{uml91CSa;4dbvbne3vzbybw-2bC:t|gl|bbxep9uI:e:F=Da/+lU0n7pS=bbTa+VEaqq8b>x,8W?384X8bSxTa9XPv,vD@;JgbWa/,7e>v9<6>y|ybfqY4h|jbW|0ojmilLzZIgbe<Nam5Cas?sGgblt/bCa+Y-bwb>w:sc*1bO-HEA"));
$write("%s",("QaItbUaeU2RN*Waj+EaT:uuunf4JtZaR<2bFaGxm,XF.bBqLp<sVa/sGyamq0n=,7v02bVaPqq5BqTaW..yV|zpN<6.6n<sVa?aBslr4qlbl5xyN*ACBa3*7*hN4Q*6@ai+3bP45OMETac+SaH:HxXlt?PaFE**6b|kgC1bVL9>\\\\{7nDMp0w|QilUk=.AyCyUkS7D;a;kbX0<a-VZa2o7zss\\\\}zGl038bv73SrhRBL\\\\{Au/glsYa\\\\{HHpsN@\\\\{1=ueO@M@\\\\}m@/|>xnk.9Y@G1w+ZM;z3.bfDV/MGOIWa-b4v6j3ptOd\\\\}@GuZ.KwZ\\\\{oR:lb*7Bowb=rvIzZ,pAq*9Rats.HXs1b4vZYz+2220PXfbNx5bZmfZhb:7Y5ibN?PhTaOao-wziXBqNIi\\\\}9L0|,1>ao/s,3z6nNa6cN*R:.b7eXFItTaWaUFVa6jg@EaS5Ol+Bx/OaA@c.r=PXvcV\\\\{.@\\\\{9OaGnnysm>np*xn3\\\\{Da0?<@\\\\}2e/zb>awlI@>*6bU,hm*\\\\{Fa?,Eajy7y2qHxf<HuauUtKXc.TaR+DsrQL1vp9*/u*bNa3>76*m8L/\\\\{0b.+c.dX@Xlb<BOILKo0A.ybN=vcPL*=PquWN01pr=.b*bhw*b\\\\}X26glxb2XLsVa+y6b.b0bwz\\\\}ttrOajmqshwgzMCo.XaybK,w\\\\{R\\\\{jbsvwyab\\\\}6XrMse3cy8bIePms?hbslRWTwY8GaMOSaLnVATogm8+wbxb"));
$write("%s",("W1D3CaQaXb|QXp,WEo?NJVu\\\\{Ed7@zl=atqFpKuLun3rQ9@sn/CdbjNLnK=,cR0Ra\\\\}qUutlcIbWdN/b*bwb>aGmy+S2Fa@uwC1U\\\\{wLutba;G1@3f1O9q/BN3buOiAsGNt+bRkal\\\\{pAVDL/b.b<l0mW\\\\{it?akNzbzlyDuUnwf7\\\\}b-b|n?\\\\}Fa34-bb6rmA.ar/R,blbKtSAHdInQavb\\\\}m31Eaky6b5z3zu50zoQkxgSzp\\\\}rrJNal5ZQ4l*nWLe8tb39sGOa6thGnV\\\\}blVeb;Ugn+MeA\\\\{b8HQsPT+b<ajT.bf+EtnUrNmbBaD0@-ebw1YaA>IJ+r:mM.<aq@lbO+GQc1(f\\\\{#cw3VaGCrN8|Lz?awBdbk?4p+MI2k?OzTaPdYwPau\\\\}tbnKD9W9kE20|OvbyJab-.Mc4b7tZaWa2J|xaulT@pQaWBCa\\\\}bgmYaqmyb*?ybb\\\\{Qa3SQDtbN<4ny4NN2;z+mnbb8yhGaPglebSHFa<uhGAr3c6c1bj/\\\\}FcyvbILe2lHxejb7esMEoV3>\\\\}\\\\}T.wWrS|uTC:@\\\\{Aa4btwOaqc37U;l>xb?ddv\\\\{bTo,ukb4bm,MK7>;y.2vbK*L71tPQmeGabAueNairT|C@l>ynDmyK186|ubWmy4fLzbBNh;/zKsPq5sfvRs+\\\\{abNFSaAaNFwbuwe<TtCqZ=En|bM:aEA@zokx6SVx763Mh80;Clhb;cmcT77emP\\\\{FSoOMx\\\\}"));
$write("%s",("DJ\\\\{bc**pq/hwky,+6cJ,\\\\}A.\"\"),\"& VbLf &\"(\"\"nF*i+6d5.,1XQZ*=@fbA.8bG\\\\{/KIltb3pD3H?*p7n.,jrPl9F,QquhycyOw9bpRwnLQwEjBX.H/+b=apBWEL1\\\\}62MX4t<\\\\}bi9Da,bpMQ\\\\}Xa5;>aj<u|628+Ga68t,2.D>G;/v9|6b?afPGAPab7OaN>PlWn\\\\{H@6ebBsGIR-TsSa>oS.1b1b6=2*S*=aebR-Ra<oty<*RaVt6=d5Ul@34b,.>.x\\\\}abxbtwA.mn6xvI<|1bnJx\\\\}fb=nmEm,.-2*2*/CboI*@|C,-r0*c</yVzY4zbU4|u,bvHwo7b\\\\{b0r3*m+Wamb4bK*4hNa*bn35;Ta.b@qkplbd,Pa/bue<umFsls\\\\{3bOtWumu@a<*r.pMWaM5-|U*u|HE22LFh+=axblbCa1b:rX11bxs9bBaJpbo+bFanl0qub\\\\{zk28+F6AuV|Da9EN1\\\\{1WJG|SaK\\\\{7bX\\\\{2v>aXAabmskbUacf\\\\{1<aibVv\\\\}m7wibA7+bM/I6700\\\\}bnybC-n@38i=-b/b23flOsk7+l\\\\}b1ui0,:2yLr72TE>alrVvvK6bxbM\\\\}YpOqi+xzWaQHTayzgspM<|Raebe2AKWaQ3SaN*Qkh+Ua1x+bS2<|c\\\\}+/4b\\\\}teb2bZdvbk4BqX7Saeb>4=sPC\\\\}lEEcNEaGA50ub?->aWa/bHGZM49N4Da07NaAMxywblrYas,gsmb"));
$write("%s",("J\\\\}Q6=aCxDaHnNa2b8b>aX|PL.bFyNaxbVaCatL\\\\{bC:UFeb/yrJ/yxvhb>py4bbnIcbX|5hU/3>fbu*tbkwfnQrV1FaF3I-2bi9*bzbEap*-MIuV\\\\{wwxbRagbhb72ymEE>aQahb9b0*dbS|QtHAq-7b=1:0L14bTa+|d,kFG6@tQtC31bfsoLso-d8tRaP0f6>t/wY7o<eb5qg@.l5-+/Dqxbxbbb+b<o*Aeb9>Xa|\\\\{0|JLPxEt|,\\\\{bP|Rh7s5shbxl=aWa>@GBFy|x/1/b7@/b63lbFreb7x>-tL2,2bBaQaLcZITaVANaP,xyVaub=shbvbvbabwbbo<Hg;Ba-b8JwC=s/1t|8+|bIyY\\\\}hb-bvp@aM:4Eo0J5c@Ca0bMzlba;U\\\\}t;<@C6q2-9u2I|3bv\\\\{G*/bZawbY11s@afv\\\\{97bZ:oB3\\\\{Yx<A-b>af\\\\{3>8bH:wbc9T+8K6KGaPfFKEnYH|bIvOGb\\\\{7es?in209<7@mb/|M||<hbUa,b6b@aI@KrKH*\\\\{SG2bdb-bg4JmQqZ/c+.Ecbcbwbk3xuB\\\\{3b|3xnBwmbE/QF>ax1V8@a,,U3\\\\},Ga\\\\{,F\\\\{x,v,F=p94IkbRo\\\\}=<F03SoMvh2XaD\\\\}PaG>oxAay/rty|.bu\\\\{NFaIypU=6F1b-mQ\\\\}8+bbybAvub=a\\\\{baCQ*70irUaFa=|M=-bH3U0qlv>?a,<uos8.bv?.1f?2\\\\{dIK:@an:UaCaS7Qtc"));
$write("%s",("bAw4\\\\{<an|vFQa@aEG;rvImI\\\\{997llfsQGN*e2CIMIfbOGmeCa+b\\\\}2?a@Gy8excb4b3bUaqIk.<F5CSalb:rqI,6Tvmbc,zbyISkgl3babme=a+bFl\\\\}8>\\\\}7b\\\\{I@\\\\{c,*F9v,IyDK:<iZjPac+c,\\\\}8im<:gl7bw=*\\\\{HpfbBap4\\\\{bhb,q\\\\{*N*Ea1l\\\\}\\\\}f./xV0lb?a\\\\}b*x72i9gxFrJC/t0p0b>G:rK1UF9rEFstdbBa.bB7Ga\\\\{GF:gxP3Pa=sWaVa*++b.bjbLsspbbq.76Dx0zhq+-y65G5z\\\\{bK+Zq=vT3tb15jb34*d34Xxfb+AHyjHFrxbjvTsAwYxNal.f\\\\}Pa<a82=/kbb2+b\\\\{.@/qyvbDasB2DTo*1Ba3beb5zeb2?tbFaPybn2Ghb06Vzzb/b5v<oxylbbb=aa+0wals,KlM1-zM|.F5\\\\{anzGpcflRw?\\\\{,/YuCalchb7e?aVam/XF*\\\\{05Vjr?WaH8kolnXaZ<cq|x5.ADx>XaVaz+q-g\\\\{0rPaGvK=2bRa7eLn8+5bQa/t3bgb,5?a8.Va6Ak,Y93.b\\\\{7\\\\{Xa*p\\\\}lm/5b6Dj42ghbFac<u\\\\{hb,z4bhb8bGahz@1Ca\\\\{qD32blrNsCv\\\\{bCaUahbZa\\\\{be>b@NaSaLx<aptmhnt\\\\}bGaw|ebE,nx+z*44020Qr\\\\{1lb,bq-HmfE0;+bi=v2r=tbxm:9zq7wWabb9bHrM7f.2b"));
$write("%s",("G-kb.b6>;9zbql>-xbQa?3inO:sBGm-sE7vb@d7bybIr\\\\}6K3P>mbd->=T@nqztj-|y/>PaQqVa@|?nl*,:n=a0iE0bgE*b*bEBaD*\\\\}vn>z?-5;NaT\\\\}e?Tar=8+9-CwYqxbeb9bubEabfEaCw,:9DQr*?m-Cw:DVwH8cbQrDmy>PrMmGaq=Mx-:hp9b4bRaCaWbYqkh=a7bH8kt\\\\}bSqLv;uQ,H?ecFa5b.b4pU:I*<a6bypFr5b-s-,T\\\\{Ys,bJs5b4>MsaClbc7rC/C57Wadlc<q@Dp,omrGpc+EBvbRaI@UaxbWkb2\\\\{bn:7y7e\\\\{;|t8bIl2b4b3y-bt\\\\}XBVdRsvCIe3s1BX:-b5hM;jn7etfUa+=Jwso3sV|;8R+spc\\\\{3/M;lbBa1==aJc|bgn0z\\\\{:*\\\\{Y10:|v8bX\\\\{8+fbX<*9GrSBQB8bncgbwbhbCsry|vyb7bG>bqqm@d7e<4tbPq3;vl3bYxfbEsfsH4jA+b8B-pao|b7?wBncUa<A5bCa0mtbGs+biw?d5q1|**NaWx4\\\\}d.+bCwS=UacbEh4\\\\{AwdbjbAmYadbFaubFwP\\\\{*pUaY/7er=DqHrmcL>V0-bN\\\\}kbQ,Ea2b<@ub|b*b7b7l,*-bYpvbCyEpTagbP4zb8b|b<|QwJw?aQ,5;OaP,Zjab,=\\\\}pTasoX=u8M7GaV*wbM=zb5tCavb2b:rYs@rm2.,xbT*kb\\\\{hvvEm1/Ix6bEa?a=@5hOa\\\\{b,"));
$write("%s",("yzp@a8+7b7e|b@,2b/1TaGaV>1|Oao=p<FaKm\\\\{hub20<uxlDoPaWv9@1sno6bOa1btb8zhbGaL=<aI6,4-bso\\\\{b<y2;+ymw>aS?5b=svbzb+ynsE\\\\{es,bc|9b3b7e\\\\}oi5aqppebPpXa74jbRadb4\\\\{db3/d>\\\\}?bbUa-|A.mzQaYa7evb76Uaj=,-xo3bf9cnR-K|7e,tO2loO24p4bhn1?gnXaBqamPqB<,+R+FnAqOr<oXav?/bnoMh1bhnebUamb5oA.Y1=9Zd7e0bp;kb>mcq-s<45b?-mb\\\\}b.bcnOwSaQaM\\\\{n3PaProeZ9s-tbTaRmu3wo8+Pm\\\\}6Z/7e@qll/gvq@-4\\\\{0bW9lbY\\\\{jbabqn\\\\{;KrUaY+r+Eabppm\\\\{by47oZa0b8tZj>u1bd+eb/b1<rr0be<z2|o7bl>CfCo-bcn@a.bHpH\\\\}v70bY0zbD/+:Hv+|5bZj4wwbBagb15?a?ng<?aq1ubGa,lPmNtZyL5>anx2xfbspEa=r+nO2+nUa7ewbRaW;ol\\\\{m4blb?3d=/bb=lb-r+rmbIl\\\\{u*mUlib<*PaSafb/*ibE.\\\\{bG;dbO9Fadb\\\\{b7b0bEneb|,+/:*@am+j2!![2aba!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"g3b[2lpa\\\\})1(f\\\\{#(tnirP;)23&Z0Da?a7e2b*b>aPa;;6|ybdbYa/oYrRaB7?\\\\}\\\\{h1bg,2bTa0lSa@aPa8+8bub?\\\\}wmXzkb3|8:F:5bT;mb5\\\\{=91b\\\\{;Oajb,z\\\\}6Cyfb2bibjlscYat<amAoSofc1<mbNaxykbdqF94b,bR|Ea-b1bAoUatlzbS|-bVa+h|\\\\{Dvmbtb,5zlam*;>a=/hb,bXa-bG;=a9bdbL76mXa2b6bvbL7mwO20fm,tfZ6wbvo7b|\\\\{D4Z|8bQaDaNaO2/,GpAq0|vp>a?n<ajbj8Kzxo\\\\}tNalbxbZaGa?l5\\\\{q/6gP\\\\{ibuby|\\\\{jZa2bA7yprq*4O2cbe;Za+bhb;5no;5Ca3b@a5xhb?afbfb;3Tt43Pa-bvbm,Va>aKqTar1lb+/pv+bktQaB1Ba8+cbTarhxb7bqtcbq14b4b\\\\}b=avvzb5bwbibWaYk3-D\\\\}9.nu-b\\\\{:5bAaDm8bab-bJ9nuMpSs0w.wr:jrY,cyVjHy@uVz4b9vzb7btwl./y-bVjebwbSa=i\\\\}yE/bb4bbb\\\\{b-bOzL9<\\\\}zbB\\\\}isD9OaYj:rl.Yjmtw2/bHbOans-bubVa7iybe2:wVa+eQa>aA0Fn:t*bdbPawbn9l9Xap*5vvbxm=amb?-+|Sa|bYan/-mvbVa<aCqZoH1+bClkb=aibfwl|YaG|Paubl*YkcbU"));
$write("%s",("aK\\\\{Ow?ayb,\\\\}1bybBm@m5o;m?\\\\{rrb\\\\{wm/qDa;7xbgbt\\\\{Z4B18+-mvtV0>aq/urvmb-jb.-\\\\}bwb|,Va@aBuibKhZaOrez/bjb?n7xzbSa/qyblsBai2*bBx<a1n*b\\\\{jJ\\\\{k|Eo@1@r8x;4+bvb,bIw6bDaD.7-Oz36O6,bhbzbibg4cbFa.bArAqGsEvYakbGnYkWkkbefzrwb\\\\}\\\\}Pa3bmbzbabdnQqhb2bbbQaalB5Qajb5,bbIxS\\\\{4b@d>17i7be*\\\\{fYa<rwbd586\\\\}by60bUuAaQvQtabO6W3W\\\\{Y\\\\{-m4bUzTaPab\\\\{5b1bubjbPaEvQa*d*1copm.babVlSaNam/eb8b5bcbR4Qq8bbbtb-matpubbww2,Da8bjbSa+w\\\\{b8+mbvbjbZawr\\\\{mgbFasmBa,bx/mbubVvEaxb7el\\\\{j\\\\{mb@2e\\\\{zbv5gbab\\\\{bHpR-wvurk1b\\\\{9bUl\\\\}mub8bxb:o>o|*1bLoFpAa>acbLrJrHr1bY+Eas+rt@aebhbmbwbCvT1+m0f+\\\\{3zX1ybntWa<acb5xGrYa|/wzD*Oz;36w<uW0TyfbmbN*bf\\\\}l1b8*efjbW.c+Jr20yb<m+b0babQte0<aabcmzb0b1bsrl*fbe2L|5s8tbb:vy01+xbEa|by2e2nxZaimXa7yZa-zjbf.sv/tzbtbAa1+Ya=m7e7eVl;4/lYsNadbkbjb3thb3,xb*b,b>aub8+jvt0"));
$write("%s",("Q1d-GqRa\\\\{f0b.bb|i4\\\\{bUadqAtmqLp7iRa:rrv,q6gOaSowbZaabUacz9sib6bimtt<\\\\}7cluplQ,yb+babRaH,WaQa=aiqy0>nHsRa@3Q*xyhbVaZaFa/bVa-bFa=ajb-b6.2b=s6bKzZa5b;r0bMm0b+rBatb82GbBz6nYoMvR-erZaBa-ycbe2jb1smedbMmnoon?aGmpeflEv.\\\\{Wy|x7yybtbBd*b3bmt\\\\{bcbN|:qCa+mXa30HvDwkb<uTaUa7bI|eb\\\\{bX\\\\{Ap.-i/GaH.i\\\\{g\\\\{.0,05bd1Bd2,PyFatbvb/boolnVaIdF/Gq8+\\\\{oF1>x|bbb|xwokbXaubtb6bybTaDm?acfabDq/y/b\\\\}b4bwbwbAa=aV/lbab>.2bYtu\\\\{kbTa7bQa/b7eubLp,b|1z1abzbjbxbH\\\\}fs,b.bXaBmY/8b+bWb-b8bBa1q/btbbzE\\\\{wbk,ZamqP|lb8rw0.bAajb*v7bjb0b\\\\}b@atb=/ucwbVa/bh,flRu*bWa1b0bgw\\\\{bIq0fNa-yeb*b\\\\{bUz\\\\}0|,fb7-?gWaNa|bkbibTt5bhbAax\\\\}0btbAx,b?x7wdtbtszQm,oNa<tcbybXt\\\\}qSal.Za/b0b5bu*bbbb.bGzcb/bab*\\\\}f\\\\{d\\\\{Wa\\\\}bUzGaSzQqKrE-,b-sVaUamu-->n?,lbDl|bi\\\\}-zbb8+Jxfbs\\\\{Kp6sybmbPxG|ib>a\\\\}b@uWw|byb/q@ae"));
$write("%s",("xfbBo<pJgWaDa5bVa<\\\\}9bUaub+b1.p*F.v\\\\{7b,bGoibDa6x|bRanqtbcy/b|bWaD\\\\}5bDaHx?fi\\\\}EaTa;u;,+bPabycb*bubAarz2\\\\}3o@-vb4q0bTajbbbf\\\\}6bPaDz\\\\}bzbdbNtB-I\\\\}2nRphbjbjb-wUa4lRaXaAa6xOaebzbQaib5bTzlbszfbFaEa5n1pYaUakt5btbfnxbAu/bmbBombgbz|hb|b>aHx@ae\\\\{mbmnCa@*S-UzgbcrFaSaSaQxgo5xU-8bOa0x4b5tOwAa.b7*4bq-Patbkxzbvb>aHdSaC*r|m+H-RaAu/y5b8+dbabgb5-to;u@-=a<uOwhx\\\\}b9bzbAa?,2bDaAas-i\\\\}xo2bAaHr7eTatb=n0bP\\\\{@rgbjnDa6btb3b9,e\\\\}DaBahbSqav1bpc6zin4bFalbtb7bbfOaOacbLlooTt7e9bZaCfYk*b1x2*7e-pTn6bZaEair-m8bDazrhb2x-btbXaFlvbOaBwOa0zRa|bOaabybfbxbAlAaYx3bAt4m6rTavbZa9bXarz2b@a>a<a+biq-d7eeb6bum|b7b=mXlZaXaPas\\\\}cbxbHpFaYalb\\\\}bY+lbYa9rEaYaRaabubPqvbspCm+n@q0boe.bDaEaGaponoEaPajb:\\\\}Aagb7ekb|m+r>+f|Zy9nTqysMr,zT*4ao\\\\}zbqt7cfn-z4bCa*bYaxb<aFa/oPazo.b3*.bBa<|VpC*@a3bZajbF*"));
$write("%s",("K*D*B*@a@*xzVaWaSaVaSa?a7blbN*SaibGa6vno=a8qlb@aTxhb\\\\{bgsRar|.bUaTa=aGd|b2b=*0tTa@t0*8b3b.bxySaWaRa?amblb/*wyWaPaWa@aSaEa=ayb6b|\\\\{Tabt\\\\{bdb>aVwYa6b\\\\}bSa=sbt5babbbhbP\\\\{Wm-bbsabRu@nXtH\\\\}>aBrmb4z:q8qybAa0fPp\\\\}bgbQa1\\\\{gbCa7bxbdb/bDrVaab4b8r\\\\}bBdab>wYajo2\\\\{ubbbEpgbgb+bYakhL\\\\{BdQfBae\\\\{?aibdbEaRawbNatbgbAaBliq8xwbFa:vBn.bxb+b\\\\}bY\\\\{Xh@zTaV\\\\{T\\\\{s|P\\\\{ab:rvqbbebRa+bn|hpAaeb5bNa0b\\\\}|jblbeb\\\\}r0bAugsvbdb0bwbebZafb+|vz4w-oUaP\\\\{DaRa*b@aUa<a<ambZa+|NaTojbtb4zkbfbtb*\\\\{mbP\\\\{|btnP\\\\{QrJpktfb7eYatbVa=auxebSa+bwbXanrTa8b|\\\\{FaRaZatbHx<aOaXa<aKtmbTa-b=aVajb=aCa/ltbgw,y3bjqYa>a.b7\\\\{6b0bYaFa,c6bzbWaBaAa|l9b1sVa8bZa=albXaQa+b@ajb6mwb-bfq\\\\}vcbEa=n/bvbNa@u0wBawbzb3bEamx>a,bYpdqzwXbzbwbrvgbNa7b4bfb\\\\{bAatwub,r*v\\\\{b5bdb7eQaBazbTaXasp6b*bUazb\\\\}bOatbHrvzxbXazbg"));
$write("%s",("kaxgbtb8b.b:rRoxb0b6bVaBaab/b+b=mibNajbwbCa5bybzbltVa:vWalbRa0b9bybXa7bhbWa1wZrcbeb<aYa-l*b<a@aDa=aGaEuoxxbPa@dTa;y@a/y8yfu2blb2bplib5vrrdbNa8b\\\\{bjb9pCqjbyb@aBa|bjbxuOa0b0y.yvbCa|bib+bGs/b@akbgbybZakbNa,b2bCa6lovUaEaEaAaWaUaAa2bXaYaWa>a0b3bxbAaDafbrmPohwabib*bSx+b>ambGamomb.bYa*vmb7eibSaXaRabbdbCwjb\\\\{by!![2aba!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"g3b[2lpa\\\\})1(f\\\\{#(tnirP;)23&=,bWoAaubgbkb?pabTaLs>s\\\\{ecbTkAaCaVa3b+plbAalbgbvbSa6bebPr*bfb7bSa@vAejtsrCaTaqs@uTtCpQabbFaebqpFa7exm3bkbVw@aQp4ack8uSa.bRacbAakb1o,bkbQaPa8b:wEvGoWrYa9bls,s*b/bXaab.bwbPvRfWaMmevqpkb*v|v7bRaKp6bYa4qubXaCadb+b1hPaBv@v>vkbkbKu4bdbrmtbdbVa7banApgo\\\\}blbTn+b6b,babXa"));
$write("%s",("4bGsye?p+l1b7ezo?adb.bSaCabbLs?a8vFrMpBacbKuvv7b.bFaTkvbPazbOaCafb6b2b-bQa-tCacbBnnopqZaQatbEanc*dDa2cJuGaCtRaubkbunYk3bSaub>tUaDmmbibumeblbwctbkhYs*b4q2bueQa8b6bUa9bPa>akbIe2bZa-bbbtq=a0buqQaMmcb\\\\{bib1bQa6b<a7eab3b1l>fwbabZaAa3bubmb4afpSrBaku<s5htlib0bVpyb?aSoUqSqpc=aabOa7eCfjbOqTs@a@awb?aXaOakt1bUawbUa/bPpBa1b\\\\}b/blbTmzrBaubWatb;q/bcbbbMg,bPaUoNacbXk\\\\}b7bcbSaJrLl+b8b7edbRqXambvr7b3b,bfb8bHq\\\\}b\\\\{b2b1bTakbSqOaWajb3lTaBa0b|bUaybjsOafbab-mfbbbZamb=a1bvbhsdb5b3bYagb|bSn<aXajm=afb4bybbo\\\\{bwbgb*b2bYaNa\\\\{blbvbXahbPa0bzbXa|b,bNavb<aCaFa8bUn<mcbBaFa*bps7eFaOaAavb*b+b,bOa,b5hFals1b,b/bEa:rjhdfCfVa+b-b@aYjAa\\\\}bfb+bybismbmbSaybcb8bypVaQa2b>a3rmbKmbb/b6b4b1rubnmdpab0b-b<aTa*bTa0bkbPa4bubPa=qBabb-bebFajokqZaMpXaZa,bSa/b>a*peb|b\\\\}bYaVa7e8b7btbtbEpWaEajrvbub4oy"));
$write("%s",("bgb3b\\\\{bzblb*bxnbblbibjbTm8b2bfb*b=aYa;pPaNaCa8bWa7bwbbpimjb7bXajbcbPa,o,b\\\\}bxb/bCfXa1b*babFaUaOa|bEacb1b7b0f8bebXaDa2bmbXacbPp9bmb7bZaVakb9bbbKp5bTaubvbjhKpkbebPoCa/bafWa5bYacbibEa1bab\\\\}babhbwb;o\"\"),\"& VbLf &\"(\"\"2bPa|b6bto?a/b<pOa>abbSlIm=a-b0b2c3b0bcb?a3bTacbmb\\\\{bbbfbUaib,bebmbUnRa5b/c9b0bubNa\\\\}bVatbfbwb\\\\{b>l3b|bTaZagb8b,bFawb.bCaOaxbDa.bkb7mjb.bTnubfbzb@ahoab1bXhVheknmkbWacbXa6b5b,bWaCaebkb|babQaTa\\\\{bao?axmFamlEaebTaQa1bfbOa8bgljhRavn@a/bPa?amn<a,b=mub7bNaWakbzbYaXabb3b7babcb\\\\}bvbbbOa/bDakbFa|bMm7e?dub7e\\\\}bDallwbaf?a\\\\{bBaRaKl\\\\{bkbxbAe>a*lTaAd-b\\\\{bYajb9b.b?aebPalbwllbwbybkbZa4bDa\\\\{jibIdPa,bwbkbynwnunlb6g2b0bQaybLmGaTeEaOa6b9b4mRaPadb7b/b5bOaYa0b7bVaXa+bOa\\\\}bXm<aUa3bPaibTadbmbhbTa\\\\}b:mXa>aUa\\\\}bUaRm@awlub\\\\{bUd|bDaUaPa7bDa@aFa1bWaql7bbbYaa"));
$write("%s",("bvb@aYaEa,b0bZa\\\\}b0bWa1lvb6bNaDazb=a>axbhb*bXaEaDaFa3bjb>azbDaDa3bAa0bdbDa|bAaFaQa4almdkfk9btbbb|bhbDajbQa?a,bZahbhb4bEadbib/l-l+l+dkbdbLcbbablbmb>agbBa5b>awb6bmb*b7e7b<a>adbdbefYa4l|b4bxbybPaGijbTaab@a7e1bebgbjb,b-b6b+hebQa7eql,bTa>aFajb\\\\{c>a7bdbCaEaybVdQa4bSa>aDa*bibBadb9b*b-bEa7b6bAaEaKk.kSi6ipkkkAkGi-a+jNj5kZhai/k9kFdQilk1k;afiykskRioj.jYiwk6iuk\\\\}kzjLjxkdjCaCeMjjkwbXbNi>jRjliji@jSj8jEajitj-iHiFi3j?jKj@i4aWhbk9aXhHfUh/b-b4bCeEfub+eNi+jEj7jbjdhAj-jZd=jhi9aEa.i9jxj0j-ahg4jDi,juh*jwd:azjlj1j=aAaojuj3iyjejkiajPimjPaxhkj<g<a-bfiMirjjjaj5iOifj9i+ibjMfZiNidhLicj:aCaaiCiTi>aAa-a*f|iIi+i9aai:i,iAaEdxfEigi2ihgBizbmizi8iBaCe4iuiIh0i*bNcsf-d5bxbfi1inixi@axfii\\\\{b\\\\{ipi*fsiOaaitiyi?aAaxfviaieimiFajihifioidi9afiHaSeSh8aCa@aCe1b+d8aZhMe8arb8a8a2b4a4a3aGf4a-exb3bHb"));
$write("%s",("6bxfCgzbxbubHaMfFgreIg3b4b.b-e,cCe\\\\{c1bzb.b1b\\\\{h/hvhthNg?a=aGf8btbhhthKfRgzg>aBamgYf?atg+gOb\\\\}gZdobfhogBa?amg|b|bvbaf.b3b>bTdObchTe*g\\\\{gcgEdmgzbIbEfrb3bzejgegrgMfpg@aCamg2b3btf:b*f7fSeQeIb:cCewd-b3a?a@a3aKa\\\\{b;apcwbxeIa3b1b?f,b|b0aTdZcWeSbgghgsgHf@aagBe@eTdYcJffg*fdgBaGf-eybYfXeNf5fLfreSeIfDa3a3fifOe1aEc1aSbRbubwb7e,btePa/eUe*fRe3a>a3a1bxewb+bxfPefc/b8b1bJbxb;a:bSesdZdEc.eSe<e;cZaxfrffc5baeVewfoctbxe-aSeNd6c4c/bCewbAe3b|c;a<bre:bre3bCe8b5c,bxb2b2btb;a?aie:eZc8ePa9e3e-eJbvdHareKe6dGa6exb-b6c4a-are.b\\\\{bmcMajare-breZddd2eGa+b-dtereGa5aZdYc?cre4c2bzb;azb-bHb3b2bJa7b?aSdaeYdRaYaOaVafbVaibTdddRdPd-a?a;a>a-aPaBaedVaNaUa?a?aed-aebcbkdvbpbEabc7bFaAaAa?a>anb-dub.b+bzb>bMa/a?c9ajc<bFaFa9a>a:b;ajcIc+b+btb\\\\{bvb3b:c>bYbWbjcKbIbGb;akd6a6ajcfdedXcadDcddCbbd6a/aZcd"));
$write("%s",("dZcCcWcCcYcEcjc9a2b5aOcMcKcIcxbvbtb+b/bxb1b5a1a/aEcSb/aObic9aCbNb:aIaIbtb,b:avb|b+bub4bcb-bpcnclcHaebdbJaGaxb,btb-b8a1bxbwbtbxbUa-b.b|b3bvbxbfb/aSbnb5aIb.b\\\\}b-aIb-avb-a1b.bybHa6aCbObsb*bCbobBbNaHa3b-b|b1b/bJaNa/aob5a/a5aJa2bg[~ia3(f\\\\{#,43.3\\\\}ia9541(f\\\\{#X3~ma(f\\\\{#(tnirP;)23\\\\}ja7362(f\\\\{# [4Lma5904(f\\\\{#q\\\\})6j3bh4Tg5Mda132g7Tja5683(f\\\\{#&[2iha=s,y=z,s6[\\\\{8Qea0603+:Vba0-;\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'i6[Y3+|8jk5[-;Hba76?Uca560<a7>[u8[6=iyay,]99999[gnirtS wen=][c n3aea\\\\{)v]y3b&a(niam diov citats cilbup\\\\{RQ ssalc[4Lba7@DVea9493$?[h9Uba3~@Wba3~@bj:[9a& cdln&&&&;maertStnirP/oi/avajL tuo/metsyS/gnal/avaja:b&ategn&&&&2 kcats timil.n&&&&]; V);=:a;3ecaL[I:aD:hha dohtem;3a/4nga repus~3acaRQ83cgassalc.|>[\\\\{:Rba5>E(\\\\}9-ca14#:(i6[\\\\{:.oa(=:s;0=:c=:i;)o9ajaerudecorp>=Mba0"));
$write("%s",("$Ma>=Qba9-R[PF[g5Qca75.RUza1251(f\\\\{#&(tnirp.biL.oken\\\\{,9bianoitcnuf/G[96[A8[.3cba1BNWK;[qa(rtStup=niam\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'tni[>Nx8dkawohsn\\\\})840h;\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'MJ+ba8~7Uda332Z4Qea1918c@Xha=q\\\\})486h6Uca148GQba7f9bta(amirpmi oicDAx\\\\})42QIaca3Cl3fpani;RQ omtirogla?9Ml4bk6aea.tmf>Acfacnuf;t4Tdatmf[3Ugaropmi;|Jafagakcay>Mda115)6dbapu6Mc4bba-X3Sjatnirp tesu=MyIaca(n)BQca725:a#a,s(llAetirW;)(resUtxeTtuptuO=:$5Mca36)6ea4RdaS CZ3M.3aca&(X4Rba [5[[5SiaRQ margof5O.3ajaS D : ; Rm5Tba\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'X3Sqa. EPYT B C : ; Aj5Tka)*,*(ETIRWt5UhaA B : ;e4Sba [2cj5Vba:a4(+3[+3wda(nfKC&;Ya|a(etirwf:oin\\\\})8(f\\\\{#>-)_(niamp3cpD~ka(f\\\\{# cnirpP@~T4ahastup.OIVO,FLataM diov\\\\{noitacilppA:$[cea[06xE3k75a*Mcpadiov;oidts.dts 5Ka14\\\\{kaenil-etirw45lva(,\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'s%\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\'(gol.elosnoc;)\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\'K3s[2cya\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\' nioj.)1+n(yarrA>-)n(=ff4kia!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\}54,1\\\\{.n3cja# qes-er(YRdba&l5rba!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"$Sk$3lo3r33tla1% ecalper.S4l(3cs=gsarts(# pam(]YALPSIDq6cua!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\".NOISIVID ERUDECORPU3kma.RQ .DI-MARG~3oE3dnaNOITACIFITNEDG9dsa[tac-yzal(s[qesod(n6apa!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\");\\\\}\\\\}!\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\");\\\\}/****/e3a\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"),s[99999],*q=s;int main()\\\\{int n,m;for(;*p;)\\\\{n=(*p-5)%92+(p[1]-5)%92*87;p+=2;if(n>3999)for(m=(*p++-5)%92+6;m--;q++)*q=q[4000-n];else for(;n--;)*q++=*p++;\\\\}puts(s);return 0;\\\\}\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\");gsub(/!/,\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\",s);for(print\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"define void f(n)\\\\{\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"00g,\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";for(m=1;m<256;m*=2)\\\\"));
$write("%s",("{\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"00g,4,:\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";if(n/m%2)\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"4+\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\",\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";\\\\};\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"4,:,\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\}\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"389**6+44*6+00p45*,\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";++j<=length(s);print\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"f(\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"n\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\");\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\")for(n=9;substr(s,j,1)!=sprintf(\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"%c\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\""));
$write("%s",("\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\",++n););s=\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"4,:,\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";split(\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"145 160 17 17 17 23 252 141 0 46 125 231 229 231 250 151 243 243 243 231 231 207 159 63 4 231 249 255 191 225 17 127 206 103 51 57 152 37 255 57 204 230 103 48 79 159 159 151 252 231 51 51 57 193 47 249 204 230 102 115 4 251 190 249 243 207 57 206 115 158 9 231 57 156 206 102 9 193 48 96 "));
$write("%s",("22 236\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\",a);for(i in a)\\\\{s=s 0;for(c=a[i]+0;c;c--)s=s\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"1+\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";s=s\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\",\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";\\\\}print s\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"@\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\"));
$write("%s",("\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\nquit\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\}\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\")');\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\";FORiTO UPBtDO INTn:=ABSt[i];print(REPR(50+n%64)+c+REPR(50+n%8MOD8)+c+REPR(50+nMOD8)+b+\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"J\\\\\\\\\\\\\\\\\\\\\\\\\\\"\"\\\\\\\\\\\"\"+a)OD\\\\\\\\\\\"\"\\\\\\\\\\\"\"\\\\\\\\\\\"\");end;\\\"\")\\nsys.exit 0}\"\")]]></xsl:template></xsl:stylesheet>\":s=\"   \":For i=0To 7:s &=Chr(32-(Asc(c)>>7-i And 1)*23):Next:System.Console.Write(s &n &Chr(9)&n &\"  \"):Next:System.Console.Write(n &n &n):End Sub:End Module"));
end endmodule